* NGSPICE file created from wrapped_snn.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

.subckt wrapped_snn active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vccd1 vssd1 wb_clk_i
XFILLER_79_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09671_ _15674_/Q _09679_/C _09583_/X vssd1 vssd1 vccd1 vccd1 _09674_/B sky130_fd_sc_hd__a21o_1
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08622_ _08622_/A _08622_/B vssd1 vssd1 vccd1 vccd1 _08623_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08553_ _10697_/A vssd1 vssd1 vccd1 vccd1 _08554_/A sky130_fd_sc_hd__buf_2
X_08484_ _08484_/A vssd1 vssd1 vccd1 vccd1 _08485_/B sky130_fd_sc_hd__inv_2
X_09105_ _15559_/Q _09145_/B _09110_/C vssd1 vssd1 vccd1 vccd1 _09112_/A sky130_fd_sc_hd__and3_1
XFILLER_109_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ _08872_/X _09029_/B _09032_/B _09035_/Y vssd1 vssd1 vccd1 vccd1 _15539_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_89_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09938_ _09938_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _15722_/D sky130_fd_sc_hd__nor2_1
X_09869_ _09869_/A _09869_/B _09869_/C vssd1 vssd1 vccd1 vccd1 _09870_/C sky130_fd_sc_hd__nand3_1
XFILLER_85_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11900_ _11900_/A _11900_/B vssd1 vssd1 vccd1 vccd1 _11905_/C sky130_fd_sc_hd__nor2_1
XFILLER_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12880_ _16176_/Q _12889_/C _12879_/X vssd1 vssd1 vccd1 vccd1 _12883_/B sky130_fd_sc_hd__a21o_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11829_/Y _11824_/C _11826_/Y _11827_/X vssd1 vssd1 vccd1 vccd1 _11832_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14550_ _14550_/A _14550_/B vssd1 vssd1 vccd1 vccd1 _14555_/C sky130_fd_sc_hd__nor2_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _16018_/Q _11764_/C _11591_/X vssd1 vssd1 vccd1 vccd1 _11762_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _16264_/Q _13731_/B _13507_/C vssd1 vssd1 vccd1 vccd1 _13503_/C sky130_fd_sc_hd__nand3_1
X_10713_ _10708_/B _10711_/B _08705_/B vssd1 vssd1 vccd1 vccd1 _10714_/B sky130_fd_sc_hd__o21a_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _16403_/Q _14598_/B _14486_/C vssd1 vssd1 vccd1 vccd1 _14481_/Y sky130_fd_sc_hd__nand3_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11693_/A _11693_/B _11693_/C vssd1 vssd1 vccd1 vccd1 _11694_/C sky130_fd_sc_hd__nand3_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16237_/CLK _16220_/D vssd1 vssd1 vccd1 vccd1 _16220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13432_ _13432_/A _13432_/B _13432_/C vssd1 vssd1 vccd1 vccd1 _13433_/C sky130_fd_sc_hd__or3_1
X_10644_ _15855_/Q _10652_/C _09683_/A vssd1 vssd1 vccd1 vccd1 _10644_/Y sky130_fd_sc_hd__a21oi_1
X_16151_ _16261_/CLK _16151_/D vssd1 vssd1 vccd1 vccd1 _16151_/Q sky130_fd_sc_hd__dfxtp_1
X_10575_ _10418_/X _10573_/B _10473_/X vssd1 vssd1 vccd1 vccd1 _10575_/Y sky130_fd_sc_hd__a21oi_1
X_13363_ _16245_/Q _13364_/C _13140_/X vssd1 vssd1 vccd1 vccd1 _13365_/A sky130_fd_sc_hd__a21oi_1
XFILLER_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15102_ _16503_/Q _15109_/C _08747_/A vssd1 vssd1 vccd1 vccd1 _15102_/Y sky130_fd_sc_hd__a21oi_1
X_12314_ _12371_/A _12314_/B _12320_/A vssd1 vssd1 vccd1 vccd1 _16094_/D sky130_fd_sc_hd__nor3_1
X_16082_ _16118_/CLK _16082_/D vssd1 vssd1 vccd1 vccd1 _16082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13294_ _13292_/Y _13286_/C _13290_/Y _13291_/X vssd1 vssd1 vccd1 vccd1 _13295_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15033_ _16492_/Q _15033_/B _15035_/C vssd1 vssd1 vccd1 vccd1 _15033_/X sky130_fd_sc_hd__and3_1
XFILLER_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12245_ _12245_/A vssd1 vssd1 vccd1 vccd1 _16085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12176_ _12174_/Y _12170_/C _12172_/Y _12181_/A vssd1 vssd1 vccd1 vccd1 _12181_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ _11978_/A vssd1 vssd1 vccd1 vccd1 _11353_/B sky130_fd_sc_hd__buf_2
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15935_ _15365_/A _15935_/D vssd1 vssd1 vccd1 vccd1 _15935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11058_ _11078_/C vssd1 vssd1 vccd1 vccd1 _11093_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10009_ _15740_/Q _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10009_/X sky130_fd_sc_hd__and3_1
XFILLER_37_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15866_ _16570_/CLK _15866_/D vssd1 vssd1 vccd1 vccd1 _15866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14817_ _14813_/Y _14815_/X _14816_/Y _14811_/C vssd1 vssd1 vccd1 vccd1 _14819_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15797_ _16595_/CLK _15797_/D vssd1 vssd1 vccd1 vccd1 _15797_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14748_ _16447_/Q _14748_/B _14750_/C vssd1 vssd1 vccd1 vccd1 _14748_/X sky130_fd_sc_hd__and3_1
XFILLER_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14679_ _16435_/Q _14716_/C _14621_/X vssd1 vssd1 vccd1 vccd1 _14681_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16418_ _16595_/CLK _16418_/D vssd1 vssd1 vccd1 vccd1 _16418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16349_ _16389_/CLK _16349_/D vssd1 vssd1 vccd1 vccd1 _16349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07984_ _14000_/A _08183_/B vssd1 vssd1 vccd1 vccd1 _07986_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09723_ _09810_/A _09723_/B _09723_/C vssd1 vssd1 vccd1 vccd1 _09724_/A sky130_fd_sc_hd__and3_1
XFILLER_86_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09654_ _09647_/Y _09648_/X _09650_/B vssd1 vssd1 vccd1 vccd1 _09655_/B sky130_fd_sc_hd__o21a_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08605_ _15460_/Q _08619_/C _08604_/X vssd1 vssd1 vccd1 vccd1 _08605_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09585_ _15656_/Q _09585_/B _09592_/C vssd1 vssd1 vccd1 vccd1 _09587_/C sky130_fd_sc_hd__nand3_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08536_ _08515_/A _08515_/B _08535_/Y vssd1 vssd1 vccd1 vccd1 _08543_/A sky130_fd_sc_hd__a21o_2
XFILLER_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08467_ _08502_/A _08467_/B vssd1 vssd1 vccd1 vccd1 _08496_/B sky130_fd_sc_hd__and2_2
XFILLER_11_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08398_ _08463_/A _08463_/B vssd1 vssd1 vccd1 vccd1 _08399_/B sky130_fd_sc_hd__xor2_4
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10360_ _10755_/B vssd1 vssd1 vccd1 vccd1 _10360_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09019_ _09142_/A _09019_/B _09019_/C vssd1 vssd1 vccd1 vccd1 _09020_/A sky130_fd_sc_hd__and3_1
XFILLER_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10291_ _10338_/A _10291_/B _10291_/C vssd1 vssd1 vccd1 vccd1 _10292_/A sky130_fd_sc_hd__and3_1
XFILLER_128_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12030_ _16056_/Q _12038_/C _12029_/X vssd1 vssd1 vccd1 vccd1 _12033_/B sky130_fd_sc_hd__a21o_1
XFILLER_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13981_ _16332_/Q _14148_/B _13981_/C vssd1 vssd1 vccd1 vccd1 _13991_/A sky130_fd_sc_hd__and3_1
X_15720_ _15812_/CLK _15720_/D vssd1 vssd1 vccd1 vccd1 _15720_/Q sky130_fd_sc_hd__dfxtp_1
X_12932_ _12932_/A vssd1 vssd1 vccd1 vccd1 _14060_/A sky130_fd_sc_hd__buf_6
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16642__47 vssd1 vssd1 vccd1 vccd1 _16642__47/HI _16718_/A sky130_fd_sc_hd__conb_1
X_15651_ _15791_/CLK _15651_/D vssd1 vssd1 vccd1 vccd1 _15651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12863_ _12863_/A _12863_/B vssd1 vssd1 vccd1 vccd1 _12868_/C sky130_fd_sc_hd__nor2_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _16423_/Q _14603_/C _14544_/X vssd1 vssd1 vccd1 vccd1 _14604_/A sky130_fd_sc_hd__a21oi_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11814_ _16025_/Q _11922_/B _11814_/C vssd1 vssd1 vccd1 vccd1 _11814_/X sky130_fd_sc_hd__and3_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _16551_/CLK _15582_/D vssd1 vssd1 vccd1 vccd1 _15582_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12790_/Y _12800_/A _12793_/Y _12788_/C vssd1 vssd1 vccd1 vccd1 _12796_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14529_/Y _14531_/X _14532_/Y _14527_/C vssd1 vssd1 vccd1 vccd1 _14535_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _12312_/A vssd1 vssd1 vccd1 vccd1 _11969_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464_ _16402_/Q _14464_/B _14466_/C vssd1 vssd1 vccd1 vccd1 _14464_/X sky130_fd_sc_hd__and3_1
X_11676_ _11957_/A vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16203_ _16237_/CLK _16203_/D vssd1 vssd1 vccd1 vccd1 _16203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13415_ _16252_/Q _13424_/C _13414_/X vssd1 vssd1 vccd1 vccd1 _13415_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10627_ _10639_/C vssd1 vssd1 vccd1 vccd1 _10652_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14395_ _14427_/C vssd1 vssd1 vccd1 vccd1 _14433_/C sky130_fd_sc_hd__clkbuf_2
X_16134_ _16555_/Q _16134_/D vssd1 vssd1 vccd1 vccd1 _16134_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13346_ _13344_/Y _13339_/C _13341_/Y _13342_/X vssd1 vssd1 vccd1 vccd1 _13347_/C
+ sky130_fd_sc_hd__a211o_1
X_10558_ _15838_/Q _10565_/C _10454_/X vssd1 vssd1 vccd1 vccd1 _10558_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16065_ _16118_/CLK _16065_/D vssd1 vssd1 vccd1 vccd1 _16065_/Q sky130_fd_sc_hd__dfxtp_1
X_13277_ _16232_/Q _13445_/B _13283_/C vssd1 vssd1 vccd1 vccd1 _13279_/C sky130_fd_sc_hd__nand3_1
X_10489_ _10489_/A _10489_/B _10489_/C vssd1 vssd1 vccd1 vccd1 _10490_/C sky130_fd_sc_hd__nand3_1
X_15016_ _15049_/C vssd1 vssd1 vccd1 vccd1 _15055_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_142_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12228_ _12224_/Y _12234_/A _12227_/Y _12222_/C vssd1 vssd1 vccd1 vccd1 _12230_/B
+ sky130_fd_sc_hd__o211a_1
X_12159_ _16074_/Q _12210_/B _12160_/C vssd1 vssd1 vccd1 vccd1 _12159_/X sky130_fd_sc_hd__and3_1
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15918_ _15365_/A _15918_/D vssd1 vssd1 vccd1 vccd1 _15918_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15849_ _16595_/CLK _15849_/D vssd1 vssd1 vccd1 vccd1 _15849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09370_ _15612_/Q _09371_/C _09369_/X vssd1 vssd1 vccd1 vccd1 _09370_/Y sky130_fd_sc_hd__a21oi_1
X_08321_ _08321_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08321_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08252_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__nor2_2
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08183_ _14000_/A _08183_/B vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__or2_1
XFILLER_146_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07967_ _16578_/Q _08178_/B vssd1 vssd1 vccd1 vccd1 _07968_/B sky130_fd_sc_hd__xnor2_4
XFILLER_114_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09706_ _09792_/A vssd1 vssd1 vccd1 vccd1 _09706_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07898_ _11339_/A _07898_/B vssd1 vssd1 vccd1 vccd1 _08296_/B sky130_fd_sc_hd__xnor2_1
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09637_ _09635_/Y _09642_/A _09632_/C _09633_/C vssd1 vssd1 vccd1 vccd1 _09639_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ _09656_/A _09568_/B vssd1 vssd1 vccd1 vccd1 _09568_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08519_ _08518_/Y _08428_/X _08479_/B vssd1 vssd1 vccd1 vccd1 _08519_/X sky130_fd_sc_hd__o21ba_1
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09499_ _15638_/Q _09585_/B _09507_/C vssd1 vssd1 vccd1 vccd1 _09501_/C sky130_fd_sc_hd__nand3_1
X_11530_ _11528_/Y _11529_/X _11525_/C _11526_/C vssd1 vssd1 vccd1 vccd1 _11532_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11461_ _15975_/Q _11688_/B _11473_/C vssd1 vssd1 vccd1 vccd1 _11467_/A sky130_fd_sc_hd__and3_1
XFILLER_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13200_ _13200_/A _13209_/B vssd1 vssd1 vccd1 vccd1 _13202_/A sky130_fd_sc_hd__or2_1
X_10412_ _10521_/A _10412_/B vssd1 vssd1 vccd1 vccd1 _10412_/X sky130_fd_sc_hd__or2_1
XFILLER_136_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11392_ _11431_/A _11392_/B _11392_/C vssd1 vssd1 vccd1 vccd1 _11393_/A sky130_fd_sc_hd__and3_1
XFILLER_99_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14180_ _14178_/Y _14179_/X _14175_/C _14176_/C vssd1 vssd1 vccd1 vccd1 _14182_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _13131_/A _13131_/B _13131_/C vssd1 vssd1 vccd1 vccd1 _13132_/A sky130_fd_sc_hd__and3_1
X_10343_ _10341_/Y _10342_/X _10337_/C _10338_/C vssd1 vssd1 vccd1 vccd1 _10345_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_109_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10274_ _10322_/A _10274_/B vssd1 vssd1 vccd1 vccd1 _10274_/Y sky130_fd_sc_hd__nor2_1
X_13062_ _16201_/Q _13292_/B _13062_/C vssd1 vssd1 vccd1 vccd1 _13062_/Y sky130_fd_sc_hd__nand3_1
XFILLER_124_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12013_ _12013_/A _12013_/B vssd1 vssd1 vccd1 vccd1 _12018_/C sky130_fd_sc_hd__nor2_1
XFILLER_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16752_ _16752_/A _07770_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
X_13964_ _14806_/A vssd1 vssd1 vccd1 vccd1 _14185_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _15812_/CLK _15703_/D vssd1 vssd1 vccd1 vccd1 _15703_/Q sky130_fd_sc_hd__dfxtp_1
X_12915_ _16181_/Q _12916_/C _12857_/X vssd1 vssd1 vccd1 vccd1 _12917_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13895_ _13896_/B _13896_/C _13896_/A vssd1 vssd1 vccd1 vccd1 _13897_/B sky130_fd_sc_hd__a21o_1
XFILLER_62_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15634_ _15791_/CLK _15634_/D vssd1 vssd1 vccd1 vccd1 _15634_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _12844_/Y _12839_/C _12841_/Y _12843_/X vssd1 vssd1 vccd1 vccd1 _12847_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _15812_/CLK _15565_/D vssd1 vssd1 vccd1 vccd1 _15565_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12777_/A vssd1 vssd1 vccd1 vccd1 _13009_/B sky130_fd_sc_hd__buf_2
XFILLER_42_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _16410_/Q _14742_/B _14516_/C vssd1 vssd1 vccd1 vccd1 _14516_/X sky130_fd_sc_hd__and3_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _12009_/A vssd1 vssd1 vccd1 vccd1 _11950_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15496_ _16551_/CLK _15496_/D vssd1 vssd1 vccd1 vccd1 _15496_/Q sky130_fd_sc_hd__dfxtp_1
X_14447_ _14480_/C vssd1 vssd1 vccd1 vccd1 _14486_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_30_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11659_ _11659_/A vssd1 vssd1 vccd1 vccd1 _16002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14378_ _14484_/A _14378_/B _14382_/B vssd1 vssd1 vccd1 vccd1 _16387_/D sky130_fd_sc_hd__nor3_1
XFILLER_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16117_ _16554_/Q _16117_/D vssd1 vssd1 vccd1 vccd1 _16117_/Q sky130_fd_sc_hd__dfxtp_1
X_13329_ _16240_/Q _13336_/C _13162_/X vssd1 vssd1 vccd1 vccd1 _13332_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16048_ _16118_/CLK _16048_/D vssd1 vssd1 vccd1 vccd1 _16048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08870_ _08870_/A _08870_/B vssd1 vssd1 vccd1 vccd1 _08870_/X sky130_fd_sc_hd__or2_1
XFILLER_97_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07821_ _07824_/A vssd1 vssd1 vccd1 vccd1 _07821_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09422_ _09422_/A _09422_/B vssd1 vssd1 vccd1 vccd1 _09422_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ _09749_/A _10526_/A _09347_/B _08554_/A vssd1 vssd1 vccd1 vccd1 _09354_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08304_ _15069_/A _08104_/B _08303_/X vssd1 vssd1 vccd1 vccd1 _08314_/B sky130_fd_sc_hd__o21ai_2
X_09284_ _10797_/B vssd1 vssd1 vccd1 vccd1 _15262_/B sky130_fd_sc_hd__buf_4
XFILLER_138_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08235_ _10029_/C _08047_/B _08046_/A vssd1 vssd1 vccd1 vccd1 _08237_/B sky130_fd_sc_hd__o21a_1
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08166_ _08351_/A _08165_/Y vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__or2b_1
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08097_ _15624_/Q _08288_/B vssd1 vssd1 vccd1 vccd1 _08098_/B sky130_fd_sc_hd__xnor2_2
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08999_ _08872_/X _08992_/B _08995_/B _08998_/Y vssd1 vssd1 vccd1 vccd1 _15530_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10961_ _10961_/A vssd1 vssd1 vccd1 vccd1 _15903_/D sky130_fd_sc_hd__clkbuf_1
X_12700_ _12701_/B _12701_/C _12699_/X vssd1 vssd1 vccd1 vccd1 _12702_/B sky130_fd_sc_hd__o21ai_1
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ _13680_/A vssd1 vssd1 vccd1 vccd1 _16288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10892_ _10928_/C vssd1 vssd1 vccd1 vccd1 _10934_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ _12629_/Y _12625_/C _12627_/Y _12636_/A vssd1 vssd1 vccd1 vccd1 _12636_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15350_ _15350_/A _15350_/B vssd1 vssd1 vccd1 vccd1 _15350_/X sky130_fd_sc_hd__or2_1
X_12562_ _16130_/Q _12622_/B _12569_/C vssd1 vssd1 vccd1 vccd1 _12562_/Y sky130_fd_sc_hd__nand3_1
X_14301_ _16378_/Q _14303_/C _14132_/X vssd1 vssd1 vccd1 vccd1 _14301_/Y sky130_fd_sc_hd__a21oi_1
X_11513_ _11529_/C vssd1 vssd1 vccd1 vccd1 _11536_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15281_ _15282_/A _16702_/A _15282_/C vssd1 vssd1 vccd1 vccd1 _15283_/B sky130_fd_sc_hd__o21a_1
XFILLER_129_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12493_ _16122_/Q _12493_/B _12495_/C vssd1 vssd1 vccd1 vccd1 _12493_/X sky130_fd_sc_hd__and3_1
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14232_ _14232_/A _14232_/B _14232_/C vssd1 vssd1 vccd1 vccd1 _14233_/C sky130_fd_sc_hd__nand3_1
X_11444_ _15973_/Q _11668_/B _11444_/C vssd1 vssd1 vccd1 vccd1 _11452_/B sky130_fd_sc_hd__and3_1
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _14197_/A _14163_/B _14163_/C vssd1 vssd1 vccd1 vccd1 _14164_/A sky130_fd_sc_hd__and3_1
X_11375_ _15964_/Q _11607_/B _11375_/C vssd1 vssd1 vccd1 vccd1 _11383_/A sky130_fd_sc_hd__and3_1
XFILLER_109_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13114_ _13107_/C _13108_/C _13110_/Y _13112_/X vssd1 vssd1 vccd1 vccd1 _13115_/C
+ sky130_fd_sc_hd__a211o_1
X_10326_ _15785_/Q _15784_/Q _15783_/Q _10227_/X vssd1 vssd1 vccd1 vccd1 _15795_/D
+ sky130_fd_sc_hd__o31a_1
X_14094_ _16348_/Q _14148_/B _14094_/C vssd1 vssd1 vccd1 vccd1 _14103_/A sky130_fd_sc_hd__and3_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13080_/A _13045_/B _13049_/A vssd1 vssd1 vccd1 vccd1 _16198_/D sky130_fd_sc_hd__nor3_1
XFILLER_140_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10257_ _10255_/Y _10250_/C _10253_/Y _10254_/X vssd1 vssd1 vccd1 vccd1 _10258_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10188_ _10188_/A vssd1 vssd1 vccd1 vccd1 _15770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14996_ _16484_/Q _15156_/B _15001_/C vssd1 vssd1 vccd1 vccd1 _14996_/Y sky130_fd_sc_hd__nand3_1
XFILLER_94_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16735_ _16735_/A _07841_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13947_ _16327_/Q _13989_/C _13781_/X vssd1 vssd1 vccd1 vccd1 _13949_/B sky130_fd_sc_hd__a21oi_1
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13878_ _13878_/A _13878_/B vssd1 vssd1 vccd1 vccd1 _13883_/C sky130_fd_sc_hd__nor2_1
X_15617_ _15791_/CLK _15617_/D vssd1 vssd1 vccd1 vccd1 _15617_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12829_ _12826_/Y _12828_/X _12823_/C _12824_/C vssd1 vssd1 vccd1 vccd1 _12831_/B
+ sky130_fd_sc_hd__o211ai_1
X_16597_ _16607_/CLK _16597_/D vssd1 vssd1 vccd1 vccd1 _16597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15548_ _16551_/CLK _15548_/D vssd1 vssd1 vccd1 vccd1 _15548_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15479_ _16551_/CLK _15479_/D vssd1 vssd1 vccd1 vccd1 _15479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _08020_/A _08197_/A vssd1 vssd1 vccd1 vccd1 _08149_/B sky130_fd_sc_hd__xor2_4
XFILLER_135_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09971_ _09965_/Y _09966_/X _09968_/B vssd1 vssd1 vccd1 vccd1 _09972_/B sky130_fd_sc_hd__o21a_1
XFILLER_130_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08922_ _10414_/A vssd1 vssd1 vccd1 vccd1 _09125_/A sky130_fd_sc_hd__clkbuf_4
X_16678__83 vssd1 vssd1 vccd1 vccd1 _16678__83/HI _16754_/A sky130_fd_sc_hd__conb_1
XFILLER_131_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08853_ _08853_/A vssd1 vssd1 vccd1 vccd1 _15500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07804_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07804_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08784_ _08782_/A _08782_/B _08783_/X vssd1 vssd1 vccd1 vccd1 _15484_/D sky130_fd_sc_hd__a21oi_1
XFILLER_85_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _15619_/Q _09448_/B _09405_/C vssd1 vssd1 vccd1 vccd1 _09412_/A sky130_fd_sc_hd__and3_1
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09336_ _09336_/A _09336_/B vssd1 vssd1 vccd1 vccd1 _09336_/X sky130_fd_sc_hd__or2_1
X_09267_ _15594_/Q _09416_/B _09267_/C vssd1 vssd1 vccd1 vccd1 _09276_/A sky130_fd_sc_hd__and3_1
XFILLER_138_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _08218_/A _08218_/B vssd1 vssd1 vccd1 vccd1 _08372_/B sky130_fd_sc_hd__nand2_2
X_09198_ _09193_/B _09196_/B _09117_/X vssd1 vssd1 vccd1 vccd1 _09204_/C sky130_fd_sc_hd__o21a_1
XFILLER_107_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08149_ _10178_/C _08149_/B vssd1 vssd1 vccd1 vccd1 _08149_/X sky130_fd_sc_hd__or2_1
XFILLER_106_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11160_ _12009_/A vssd1 vssd1 vccd1 vccd1 _11381_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ _10109_/A _10109_/B _10110_/X vssd1 vssd1 vccd1 vccd1 _15756_/D sky130_fd_sc_hd__a21oi_1
X_11091_ input5/X vssd1 vssd1 vccd1 vccd1 _12225_/A sky130_fd_sc_hd__clkbuf_4
X_10042_ _10042_/A vssd1 vssd1 vccd1 vccd1 _15744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14850_ _14909_/A _14850_/B _14855_/A vssd1 vssd1 vccd1 vccd1 _16461_/D sky130_fd_sc_hd__nor3_1
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13801_ _13798_/Y _13799_/X _13800_/Y _13796_/C vssd1 vssd1 vccd1 vccd1 _13803_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14781_ _14819_/A _14781_/B _14781_/C vssd1 vssd1 vccd1 vccd1 _14782_/A sky130_fd_sc_hd__and3_1
XFILLER_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11993_ _11993_/A vssd1 vssd1 vccd1 vccd1 _12218_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16520_ _16595_/CLK _16520_/D vssd1 vssd1 vccd1 vccd1 _16520_/Q sky130_fd_sc_hd__dfxtp_1
X_13732_ _13733_/B _13733_/C _13733_/A vssd1 vssd1 vccd1 vccd1 _13734_/B sky130_fd_sc_hd__a21o_1
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10944_ _11169_/A _10944_/B _10944_/C vssd1 vssd1 vccd1 vccd1 _10945_/C sky130_fd_sc_hd__or3_1
XFILLER_44_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16451_ _16595_/CLK _16451_/D vssd1 vssd1 vccd1 vccd1 _16451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13663_ _13700_/C vssd1 vssd1 vccd1 vccd1 _13709_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10875_ _15893_/Q _10878_/C _10874_/X vssd1 vssd1 vccd1 vccd1 _10879_/A sky130_fd_sc_hd__a21oi_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15402_ _16109_/Q _16108_/Q _16107_/Q _15397_/X vssd1 vssd1 vccd1 vccd1 _16584_/D
+ sky130_fd_sc_hd__o31a_1
X_12614_ _16137_/Q _12726_/B _12614_/C vssd1 vssd1 vccd1 vccd1 _12614_/Y sky130_fd_sc_hd__nand3_1
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16382_ _16389_/CLK _16382_/D vssd1 vssd1 vccd1 vccd1 _16382_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13594_ _13594_/A _13594_/B vssd1 vssd1 vccd1 vccd1 _13595_/B sky130_fd_sc_hd__nor2_1
XFILLER_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15333_ _15333_/A _15333_/B _15337_/A vssd1 vssd1 vccd1 vccd1 _16544_/D sky130_fd_sc_hd__nor3_1
X_12545_ _16129_/Q _12770_/B _12545_/C vssd1 vssd1 vccd1 vccd1 _12545_/X sky130_fd_sc_hd__and3_1
XFILLER_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15264_ _15262_/Y _15258_/C _15260_/Y _15269_/A vssd1 vssd1 vccd1 vccd1 _15269_/B
+ sky130_fd_sc_hd__a211oi_1
X_12476_ _12510_/C vssd1 vssd1 vccd1 vccd1 _12516_/C sky130_fd_sc_hd__clkbuf_2
X_14215_ _14439_/A vssd1 vssd1 vccd1 vccd1 _14256_/A sky130_fd_sc_hd__clkbuf_2
X_11427_ _15971_/Q _11654_/B _11436_/C vssd1 vssd1 vccd1 vccd1 _11427_/X sky130_fd_sc_hd__and3_1
XANTENNA_5 _13886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _16518_/Q _15248_/B _15195_/C vssd1 vssd1 vccd1 vccd1 _15195_/Y sky130_fd_sc_hd__nand3_1
X_14146_ _14146_/A vssd1 vssd1 vccd1 vccd1 _16354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11358_ _15962_/Q _11361_/C _11306_/X vssd1 vssd1 vccd1 vccd1 _11358_/Y sky130_fd_sc_hd__a21oi_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _10306_/Y _10315_/A _10308_/Y _10304_/C vssd1 vssd1 vccd1 vccd1 _10311_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14077_ _16346_/Q _14079_/C _13853_/X vssd1 vssd1 vccd1 vccd1 _14077_/Y sky130_fd_sc_hd__a21oi_1
X_11289_ _11309_/C vssd1 vssd1 vccd1 vccd1 _11322_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13028_ _16197_/Q _13082_/B _13028_/C vssd1 vssd1 vccd1 vccd1 _13036_/B sky130_fd_sc_hd__and3_1
XFILLER_67_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14979_ _14979_/A vssd1 vssd1 vccd1 vccd1 _14979_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16718_ _16718_/A _07822_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
XFILLER_35_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09121_ _09240_/A _09124_/C vssd1 vssd1 vccd1 vccd1 _09123_/A sky130_fd_sc_hd__and2_1
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09052_ _15548_/Q _09070_/C _09051_/X vssd1 vssd1 vccd1 vccd1 _09054_/B sky130_fd_sc_hd__a21oi_1
XFILLER_108_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08003_ _08003_/A _08003_/B vssd1 vssd1 vccd1 vccd1 _08004_/B sky130_fd_sc_hd__nand2_2
XFILLER_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _15729_/Q _09955_/C _08604_/A vssd1 vssd1 vccd1 vccd1 _09954_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08905_ _08946_/A _08905_/B _08909_/B vssd1 vssd1 vccd1 vccd1 _15510_/D sky130_fd_sc_hd__nor3_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _15713_/Q _09884_/C _08629_/A vssd1 vssd1 vccd1 vccd1 _09886_/B sky130_fd_sc_hd__a21o_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08921_/A _08921_/B _08836_/C vssd1 vssd1 vccd1 vccd1 _08838_/A sky130_fd_sc_hd__and3_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08767_ _08768_/B _08768_/C _08768_/A vssd1 vssd1 vccd1 vccd1 _08769_/B sky130_fd_sc_hd__a21o_1
XFILLER_85_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08698_ _09117_/A vssd1 vssd1 vccd1 vccd1 _08698_/X sky130_fd_sc_hd__buf_2
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10660_ _10660_/A _10660_/B vssd1 vssd1 vccd1 vccd1 _10661_/B sky130_fd_sc_hd__nor2_1
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09319_ _15601_/Q _09340_/C _09252_/X vssd1 vssd1 vccd1 vccd1 _09321_/B sky130_fd_sc_hd__a21oi_1
X_10591_ _10740_/A vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12330_ _16098_/Q _12332_/C _12157_/X vssd1 vssd1 vccd1 vccd1 _12330_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12261_ input2/X vssd1 vssd1 vccd1 vccd1 _13392_/A sky130_fd_sc_hd__buf_4
XFILLER_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14000_ _14000_/A vssd1 vssd1 vccd1 vccd1 _14017_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11212_ _15939_/Q _11212_/B _11217_/C vssd1 vssd1 vccd1 vccd1 _11212_/Y sky130_fd_sc_hd__nand3_1
XFILLER_107_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12192_ _12212_/C vssd1 vssd1 vccd1 vccd1 _12226_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11143_ _11993_/A vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__buf_2
XFILLER_134_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15951_ _15365_/A _15951_/D vssd1 vssd1 vccd1 vccd1 _15951_/Q sky130_fd_sc_hd__dfxtp_1
X_11074_ _11074_/A vssd1 vssd1 vccd1 vccd1 _15920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10025_ _10029_/C vssd1 vssd1 vccd1 vccd1 _10038_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14902_ _14902_/A vssd1 vssd1 vccd1 vccd1 _14918_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15882_ _16553_/Q _15882_/D vssd1 vssd1 vccd1 vccd1 _15882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14833_ _14833_/A _14833_/B vssd1 vssd1 vccd1 vccd1 _14834_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14764_ _16449_/Q _14995_/B _14764_/C vssd1 vssd1 vccd1 vccd1 _14772_/A sky130_fd_sc_hd__and3_1
XFILLER_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11976_ _11976_/A vssd1 vssd1 vccd1 vccd1 _16047_/D sky130_fd_sc_hd__clkbuf_1
X_16503_ _16607_/CLK _16503_/D vssd1 vssd1 vccd1 vccd1 _16503_/Q sky130_fd_sc_hd__dfxtp_1
X_13715_ _13881_/A vssd1 vssd1 vccd1 vccd1 _13756_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10927_ _15900_/Q _10934_/C _10866_/X vssd1 vssd1 vccd1 vccd1 _10927_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14695_ _16438_/Q _14697_/C _14694_/X vssd1 vssd1 vccd1 vccd1 _14695_/Y sky130_fd_sc_hd__a21oi_1
X_16434_ _16595_/CLK _16434_/D vssd1 vssd1 vccd1 vccd1 _16434_/Q sky130_fd_sc_hd__dfxtp_2
X_13646_ _13646_/A _13656_/B vssd1 vssd1 vccd1 vccd1 _13649_/A sky130_fd_sc_hd__or2_1
XFILLER_20_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10858_ _13183_/A vssd1 vssd1 vccd1 vccd1 _11993_/A sky130_fd_sc_hd__buf_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _16389_/CLK _16365_/D vssd1 vssd1 vccd1 vccd1 _16365_/Q sky130_fd_sc_hd__dfxtp_1
X_13577_ _13577_/A vssd1 vssd1 vccd1 vccd1 _16273_/D sky130_fd_sc_hd__clkbuf_1
X_10789_ _15881_/Q _10789_/B _10791_/C vssd1 vssd1 vccd1 vccd1 _10789_/X sky130_fd_sc_hd__and3_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15316_ _15320_/A _15316_/B vssd1 vssd1 vccd1 vccd1 _15316_/Y sky130_fd_sc_hd__nand2_1
X_12528_ _12528_/A vssd1 vssd1 vccd1 vccd1 _16125_/D sky130_fd_sc_hd__clkbuf_1
X_16296_ _16533_/Q _16296_/D vssd1 vssd1 vccd1 vccd1 _16296_/Q sky130_fd_sc_hd__dfxtp_1
X_15247_ _16528_/Q _15247_/B _15248_/C vssd1 vssd1 vccd1 vccd1 _15247_/X sky130_fd_sc_hd__and3_1
X_12459_ _12457_/Y _12453_/C _12455_/Y _12464_/A vssd1 vssd1 vccd1 vccd1 _12464_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_126_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15178_ _16516_/Q _15215_/C _08843_/A vssd1 vssd1 vccd1 vccd1 _15180_/B sky130_fd_sc_hd__a21oi_1
XFILLER_98_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14129_ _14123_/C _14124_/C _14126_/Y _14127_/X vssd1 vssd1 vccd1 vccd1 _14130_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16648__53 vssd1 vssd1 vccd1 vccd1 _16648__53/HI _16724_/A sky130_fd_sc_hd__conb_1
XFILLER_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09670_ _09718_/A _09670_/B _09674_/A vssd1 vssd1 vccd1 vccd1 _15670_/D sky130_fd_sc_hd__nor3_1
XFILLER_95_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08621_ _08621_/A _08621_/B vssd1 vssd1 vccd1 vccd1 _08622_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08552_ input8/X vssd1 vssd1 vccd1 vccd1 _10697_/A sky130_fd_sc_hd__buf_2
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08483_ _15450_/Q _08490_/A _15299_/A vssd1 vssd1 vccd1 vccd1 _08484_/A sky130_fd_sc_hd__and3_1
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09104_ _15559_/Q _09110_/C _09063_/X vssd1 vssd1 vccd1 vccd1 _09104_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09035_ _09119_/A _09042_/C vssd1 vssd1 vccd1 vccd1 _09035_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09937_ _10220_/A _09706_/X _09932_/B _09707_/X vssd1 vssd1 vccd1 vccd1 _09938_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _09869_/B _09869_/C _09869_/A vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__a21o_1
XFILLER_86_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08819_ _14806_/A vssd1 vssd1 vccd1 vccd1 _10789_/B sky130_fd_sc_hd__clkbuf_2
X_09799_ _09836_/C vssd1 vssd1 vccd1 vccd1 _09845_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _11826_/Y _11827_/X _11829_/Y _11824_/C vssd1 vssd1 vccd1 vccd1 _11832_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11761_/A vssd1 vssd1 vccd1 vccd1 _16016_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13786_/A vssd1 vssd1 vccd1 vccd1 _13731_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10710_/A _10710_/B _10711_/X vssd1 vssd1 vccd1 vccd1 _15864_/D sky130_fd_sc_hd__a21oi_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14480_ _16404_/Q _14710_/B _14480_/C vssd1 vssd1 vccd1 vccd1 _14488_/A sky130_fd_sc_hd__and3_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11692_ _11693_/B _11693_/C _11693_/A vssd1 vssd1 vccd1 vccd1 _11694_/B sky130_fd_sc_hd__a21o_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13431_ _13432_/B _13432_/C _13264_/X vssd1 vssd1 vccd1 vccd1 _13433_/B sky130_fd_sc_hd__o21ai_1
X_10643_ _10643_/A vssd1 vssd1 vccd1 vccd1 _15852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16150_ _16261_/CLK _16150_/D vssd1 vssd1 vccd1 vccd1 _16150_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13362_ _13362_/A _13362_/B _13366_/B vssd1 vssd1 vccd1 vccd1 _16243_/D sky130_fd_sc_hd__nor3_1
X_10574_ _10469_/X _10566_/B _10570_/B _10573_/Y vssd1 vssd1 vccd1 vccd1 _15838_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_127_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15101_ _15101_/A vssd1 vssd1 vccd1 vccd1 _16501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12313_ _16095_/Q _12535_/B _12325_/C vssd1 vssd1 vccd1 vccd1 _12320_/A sky130_fd_sc_hd__and3_1
XFILLER_127_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16081_ _16118_/CLK _16081_/D vssd1 vssd1 vccd1 vccd1 _16081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13293_ _13290_/Y _13291_/X _13292_/Y _13286_/C vssd1 vssd1 vccd1 vccd1 _13295_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15032_ _16492_/Q _15035_/C _14979_/X vssd1 vssd1 vccd1 vccd1 _15032_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12244_ _12283_/A _12244_/B _12244_/C vssd1 vssd1 vccd1 vccd1 _12245_/A sky130_fd_sc_hd__and3_1
XFILLER_123_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12175_ _12172_/Y _12181_/A _12174_/Y _12170_/C vssd1 vssd1 vccd1 vccd1 _12177_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11126_ _15929_/Q _11137_/C _10905_/X vssd1 vssd1 vccd1 vccd1 _11126_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15934_ _15365_/A _15934_/D vssd1 vssd1 vccd1 vccd1 _15934_/Q sky130_fd_sc_hd__dfxtp_2
X_11057_ _11070_/C vssd1 vssd1 vccd1 vccd1 _11078_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10008_ _10005_/A _10004_/Y _10005_/B vssd1 vssd1 vccd1 vccd1 _10008_/Y sky130_fd_sc_hd__o21bai_1
X_15865_ _16570_/CLK _15865_/D vssd1 vssd1 vccd1 vccd1 _15865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14816_ _16456_/Q _14875_/B _14823_/C vssd1 vssd1 vccd1 vccd1 _14816_/Y sky130_fd_sc_hd__nand3_1
XFILLER_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15796_ _16595_/CLK _15796_/D vssd1 vssd1 vccd1 vccd1 _15796_/Q sky130_fd_sc_hd__dfxtp_2
X_11959_ _11960_/B _11960_/C _11850_/X vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__o21ai_1
X_14747_ _16447_/Q _14750_/C _14694_/X vssd1 vssd1 vccd1 vccd1 _14747_/Y sky130_fd_sc_hd__a21oi_1
X_14678_ _14710_/C vssd1 vssd1 vccd1 vccd1 _14716_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_60_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16417_ input11/X _16417_/D vssd1 vssd1 vccd1 vccd1 _16417_/Q sky130_fd_sc_hd__dfxtp_1
X_13629_ _13629_/A vssd1 vssd1 vccd1 vccd1 _16281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16348_ _16389_/CLK _16348_/D vssd1 vssd1 vccd1 vccd1 _16348_/Q sky130_fd_sc_hd__dfxtp_1
X_16279_ _16533_/Q _16279_/D vssd1 vssd1 vccd1 vccd1 _16279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07983_ _11964_/A _07983_/B vssd1 vssd1 vccd1 vccd1 _08183_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09722_ _09722_/A _09722_/B _09722_/C vssd1 vssd1 vccd1 vccd1 _09723_/C sky130_fd_sc_hd__nand3_1
XFILLER_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09653_ _09647_/Y _09650_/X _09652_/Y vssd1 vssd1 vccd1 vccd1 _15665_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08604_ _08604_/A vssd1 vssd1 vccd1 vccd1 _08604_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09584_ _15656_/Q _09592_/C _09583_/X vssd1 vssd1 vccd1 vccd1 _09587_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08535_ _08535_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _08535_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08466_ _08466_/A _08466_/B vssd1 vssd1 vccd1 vccd1 _08467_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08397_ _08279_/A _08279_/B _08396_/Y vssd1 vssd1 vccd1 vccd1 _08463_/B sky130_fd_sc_hd__a21oi_2
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09018_ _09018_/A _09018_/B _09018_/C vssd1 vssd1 vccd1 vccd1 _09019_/C sky130_fd_sc_hd__nand3_1
X_10290_ _10290_/A _10290_/B _10290_/C vssd1 vssd1 vccd1 vccd1 _10291_/C sky130_fd_sc_hd__nand3_1
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13980_ _16332_/Q _13989_/C _13979_/X vssd1 vssd1 vccd1 vccd1 _13980_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12931_ _12967_/C vssd1 vssd1 vccd1 vccd1 _12975_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15650_ _15812_/CLK _15650_/D vssd1 vssd1 vccd1 vccd1 _15650_/Q sky130_fd_sc_hd__dfxtp_1
X_12862_ _12862_/A _12862_/B vssd1 vssd1 vccd1 vccd1 _12863_/B sky130_fd_sc_hd__nor2_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _16025_/Q _11821_/C _11755_/X vssd1 vssd1 vccd1 vccd1 _11813_/Y sky130_fd_sc_hd__a21oi_1
X_14601_ _14624_/A _14601_/B _14605_/B vssd1 vssd1 vccd1 vccd1 _16421_/D sky130_fd_sc_hd__nor3_1
X_15581_ _16551_/CLK _15581_/D vssd1 vssd1 vccd1 vccd1 _15581_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _16163_/Q _12911_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12793_/Y sky130_fd_sc_hd__nand3_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _16411_/Q _14591_/B _14539_/C vssd1 vssd1 vccd1 vccd1 _14532_/Y sky130_fd_sc_hd__nand3_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _16015_/Q _11785_/C _11517_/X vssd1 vssd1 vccd1 vccd1 _11747_/B sky130_fd_sc_hd__a21oi_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _16402_/Q _14466_/C _14411_/X vssd1 vssd1 vccd1 vccd1 _14463_/Y sky130_fd_sc_hd__a21oi_1
X_11675_ _11673_/A _11673_/B _11674_/X vssd1 vssd1 vccd1 vccd1 _16004_/D sky130_fd_sc_hd__a21oi_1
X_16202_ _16237_/CLK _16202_/D vssd1 vssd1 vccd1 vccd1 _16202_/Q sky130_fd_sc_hd__dfxtp_1
X_13414_ _13979_/A vssd1 vssd1 vccd1 vccd1 _13414_/X sky130_fd_sc_hd__clkbuf_2
X_10626_ _10630_/C vssd1 vssd1 vccd1 vccd1 _10639_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14394_ _14414_/C vssd1 vssd1 vccd1 vccd1 _14427_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16133_ _16554_/Q _16133_/D vssd1 vssd1 vccd1 vccd1 _16133_/Q sky130_fd_sc_hd__dfxtp_1
X_13345_ _13341_/Y _13342_/X _13344_/Y _13339_/C vssd1 vssd1 vccd1 vccd1 _13347_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_139_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10557_ _10557_/A vssd1 vssd1 vccd1 vccd1 _15835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _16118_/CLK _16064_/D vssd1 vssd1 vccd1 vccd1 _16064_/Q sky130_fd_sc_hd__dfxtp_1
X_13276_ _16232_/Q _13283_/C _13162_/X vssd1 vssd1 vccd1 vccd1 _13279_/B sky130_fd_sc_hd__a21o_1
X_10488_ _10489_/B _10489_/C _10489_/A vssd1 vssd1 vccd1 vccd1 _10490_/B sky130_fd_sc_hd__a21o_1
XFILLER_142_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15015_ _15035_/C vssd1 vssd1 vccd1 vccd1 _15049_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12227_ _16083_/Q _12347_/B _12232_/C vssd1 vssd1 vccd1 vccd1 _12227_/Y sky130_fd_sc_hd__nand3_1
X_12158_ _16074_/Q _12160_/C _12157_/X vssd1 vssd1 vccd1 vccd1 _12158_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11109_ _11169_/A _11109_/B _11109_/C vssd1 vssd1 vccd1 vccd1 _11110_/C sky130_fd_sc_hd__or3_1
XFILLER_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12089_ _12089_/A _12089_/B _12089_/C vssd1 vssd1 vccd1 vccd1 _12090_/C sky130_fd_sc_hd__nand3_1
XFILLER_49_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15917_ _15365_/A _15917_/D vssd1 vssd1 vccd1 vccd1 _15917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15848_ _16551_/CLK _15848_/D vssd1 vssd1 vccd1 vccd1 _15848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15779_ _15812_/CLK _15779_/D vssd1 vssd1 vccd1 vccd1 _15779_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08320_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08411_/A sky130_fd_sc_hd__nand2_1
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08251_ _08251_/A _08251_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08252_/B sky130_fd_sc_hd__and3_1
XFILLER_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08182_ _13777_/A _07965_/B _08181_/X vssd1 vssd1 vccd1 vccd1 _08354_/A sky130_fd_sc_hd__o21ai_1
XFILLER_146_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07966_ _08181_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08178_/B sky130_fd_sc_hd__xor2_4
XFILLER_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09705_ _09615_/X _09701_/B _09572_/X vssd1 vssd1 vccd1 vccd1 _09709_/A sky130_fd_sc_hd__a21oi_1
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07897_ _09448_/C _08116_/B vssd1 vssd1 vccd1 vccd1 _07898_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09636_ _15666_/Q _09636_/B _09636_/C vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__and3_1
XFILLER_28_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09567_ _09655_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09568_/B sky130_fd_sc_hd__and2_1
XFILLER_130_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08518_ _08518_/A vssd1 vssd1 vccd1 vccd1 _08518_/Y sky130_fd_sc_hd__inv_2
X_09498_ _15638_/Q _09507_/C _09362_/X vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__a21o_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08449_ _08449_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08504_/A sky130_fd_sc_hd__nor2_1
X_11460_ _12312_/A vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10411_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10412_/B sky130_fd_sc_hd__nor2_1
XFILLER_139_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11391_ _11452_/A _11391_/B _11391_/C vssd1 vssd1 vccd1 vccd1 _11392_/C sky130_fd_sc_hd__or3_1
X_13130_ _13128_/Y _13123_/C _13125_/Y _13127_/X vssd1 vssd1 vccd1 vccd1 _13131_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10342_ _15800_/Q _10494_/B _10342_/C vssd1 vssd1 vccd1 vccd1 _10342_/X sky130_fd_sc_hd__and3_1
XFILLER_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _14186_/A vssd1 vssd1 vccd1 vccd1 _13292_/B sky130_fd_sc_hd__buf_2
X_10273_ _10268_/B _10271_/B _10164_/X vssd1 vssd1 vccd1 vccd1 _10274_/B sky130_fd_sc_hd__o21a_1
X_12012_ _12012_/A _12012_/B vssd1 vssd1 vccd1 vccd1 _12013_/B sky130_fd_sc_hd__nor2_1
XFILLER_120_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16751_ _16751_/A _07768_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13963_ _16330_/Q _13966_/C _13853_/X vssd1 vssd1 vccd1 vccd1 _13963_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15702_ _15812_/CLK _15702_/D vssd1 vssd1 vccd1 vccd1 _15702_/Q sky130_fd_sc_hd__dfxtp_1
X_12914_ _12936_/A _12914_/B _12918_/B vssd1 vssd1 vccd1 vccd1 _16179_/D sky130_fd_sc_hd__nor3_1
X_13894_ _16320_/Q _14010_/B _13900_/C vssd1 vssd1 vccd1 vccd1 _13896_/C sky130_fd_sc_hd__nand3_1
XFILLER_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15633_ _15812_/CLK _15633_/D vssd1 vssd1 vccd1 vccd1 _15633_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ _12841_/Y _12843_/X _12844_/Y _12839_/C vssd1 vssd1 vccd1 vccd1 _12847_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _16162_/Q _12776_/B _12778_/C vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__and3_1
XFILLER_15_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15564_ _15812_/CLK _15564_/D vssd1 vssd1 vccd1 vccd1 _15564_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _16013_/Q _11729_/C _11726_/X vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__a21oi_1
X_14515_ _14799_/A vssd1 vssd1 vccd1 vccd1 _14742_/B sky130_fd_sc_hd__buf_2
XFILLER_30_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15495_ _16551_/CLK _15495_/D vssd1 vssd1 vccd1 vccd1 _15495_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11658_ _11658_/A _11658_/B _11658_/C vssd1 vssd1 vccd1 vccd1 _11659_/A sky130_fd_sc_hd__and3_1
X_14446_ _14466_/C vssd1 vssd1 vccd1 vccd1 _14480_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10609_ _10607_/Y _10603_/C _10605_/Y _10614_/A vssd1 vssd1 vccd1 vccd1 _10614_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14377_ _14375_/Y _14369_/C _14372_/Y _14382_/A vssd1 vssd1 vccd1 vccd1 _14382_/B
+ sky130_fd_sc_hd__a211oi_1
X_11589_ _11604_/A _11589_/B _11589_/C vssd1 vssd1 vccd1 vccd1 _11590_/A sky130_fd_sc_hd__and3_1
XFILLER_128_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13328_ _13362_/A _13328_/B _13332_/A vssd1 vssd1 vccd1 vccd1 _16238_/D sky130_fd_sc_hd__nor3_1
X_16116_ _16554_/Q _16116_/D vssd1 vssd1 vccd1 vccd1 _16116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16047_ _16118_/CLK _16047_/D vssd1 vssd1 vccd1 vccd1 _16047_/Q sky130_fd_sc_hd__dfxtp_1
X_13259_ _13259_/A _13259_/B vssd1 vssd1 vccd1 vccd1 _13260_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07820_ _07824_/A vssd1 vssd1 vccd1 vccd1 _07820_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09421_ _15622_/Q _09837_/A _09428_/C vssd1 vssd1 vccd1 vccd1 _09423_/B sky130_fd_sc_hd__and3_1
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _09307_/X _09347_/B _09351_/X vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__a21oi_1
XFILLER_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08303_ _08849_/C _08303_/B vssd1 vssd1 vccd1 vccd1 _08303_/X sky130_fd_sc_hd__or2_1
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09283_ _14872_/A vssd1 vssd1 vccd1 vccd1 _10797_/B sky130_fd_sc_hd__buf_2
X_08234_ _09761_/C _08059_/B _08058_/A vssd1 vssd1 vccd1 vccd1 _08237_/A sky130_fd_sc_hd__o21a_2
X_08165_ _08165_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _08165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08096_ _08096_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08288_/B sky130_fd_sc_hd__xor2_2
XFILLER_106_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08998_ _09119_/A _09003_/C vssd1 vssd1 vccd1 vccd1 _08998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07949_ _07949_/A _07949_/B vssd1 vssd1 vccd1 vccd1 _07972_/A sky130_fd_sc_hd__xor2_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10960_ _10981_/A _10960_/B _10960_/C vssd1 vssd1 vccd1 vccd1 _10961_/A sky130_fd_sc_hd__and3_1
XFILLER_90_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09619_ _09619_/A _09619_/B vssd1 vssd1 vccd1 vccd1 _15659_/D sky130_fd_sc_hd__nor2_1
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10891_ _10914_/C vssd1 vssd1 vccd1 vccd1 _10928_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12630_ _12627_/Y _12636_/A _12629_/Y _12625_/C vssd1 vssd1 vccd1 vccd1 _12632_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12561_ _16131_/Q _12784_/B _12569_/C vssd1 vssd1 vccd1 vccd1 _12561_/X sky130_fd_sc_hd__and3_1
XFILLER_12_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11512_ _16569_/Q vssd1 vssd1 vccd1 vccd1 _11529_/C sky130_fd_sc_hd__inv_2
X_14300_ _14300_/A vssd1 vssd1 vccd1 vccd1 _16376_/D sky130_fd_sc_hd__clkbuf_1
X_15280_ _16705_/A vssd1 vssd1 vccd1 vccd1 _15282_/A sky130_fd_sc_hd__inv_2
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12492_ _16122_/Q _12495_/C _12440_/X vssd1 vssd1 vccd1 vccd1 _12492_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14231_ _14232_/B _14232_/C _14232_/A vssd1 vssd1 vccd1 vccd1 _14233_/B sky130_fd_sc_hd__a21o_1
X_11443_ _12009_/A vssd1 vssd1 vccd1 vccd1 _11668_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14162_ _14276_/A _14162_/B _14162_/C vssd1 vssd1 vccd1 vccd1 _14163_/C sky130_fd_sc_hd__or3_1
X_11374_ _12225_/A vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_124_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ _13110_/Y _13112_/X _13107_/C _13108_/C vssd1 vssd1 vccd1 vccd1 _13115_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_124_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10325_ _10276_/X _10322_/B _10324_/Y vssd1 vssd1 vccd1 vccd1 _15794_/D sky130_fd_sc_hd__o21a_1
XFILLER_113_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14093_ _16348_/Q _14101_/C _13979_/X vssd1 vssd1 vccd1 vccd1 _14093_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _16199_/Q _13102_/B _13053_/C vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__and3_1
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10256_ _10253_/Y _10254_/X _10255_/Y _10250_/C vssd1 vssd1 vccd1 vccd1 _10258_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_79_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10187_ _10250_/A _10187_/B _10187_/C vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__and3_1
XFILLER_121_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14995_ _16485_/Q _14995_/B _14995_/C vssd1 vssd1 vccd1 vccd1 _15003_/A sky130_fd_sc_hd__and3_1
X_16734_ _16734_/A _07840_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13946_ _13981_/C vssd1 vssd1 vccd1 vccd1 _13989_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13877_ _13877_/A _13877_/B vssd1 vssd1 vccd1 vccd1 _13878_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15616_ _15791_/CLK _15616_/D vssd1 vssd1 vccd1 vccd1 _15616_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12828_ _16169_/Q _13053_/B _12828_/C vssd1 vssd1 vccd1 vccd1 _12828_/X sky130_fd_sc_hd__and3_1
XFILLER_62_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16596_ _16607_/CLK _16596_/D vssd1 vssd1 vccd1 vccd1 _16596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15547_ _15791_/CLK _15547_/D vssd1 vssd1 vccd1 vccd1 _15547_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12792_/C vssd1 vssd1 vccd1 vccd1 _12798_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15478_ _16551_/CLK _15478_/D vssd1 vssd1 vccd1 vccd1 _15478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14429_ _14426_/Y _14435_/A _14428_/Y _14424_/C vssd1 vssd1 vccd1 vccd1 _14431_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09970_ _09965_/Y _09968_/X _09969_/Y vssd1 vssd1 vccd1 vccd1 _15728_/D sky130_fd_sc_hd__o21a_1
XFILLER_89_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08921_ _08921_/A _08921_/B _08921_/C vssd1 vssd1 vccd1 vccd1 _08926_/A sky130_fd_sc_hd__and3_1
XFILLER_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08852_ _08940_/A _08852_/B _08852_/C vssd1 vssd1 vccd1 vccd1 _08853_/A sky130_fd_sc_hd__and3_1
XFILLER_85_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07803_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07803_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08783_ _08870_/A _08783_/B vssd1 vssd1 vccd1 vccd1 _08783_/X sky130_fd_sc_hd__or2_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09404_ _15619_/Q _09428_/C _09252_/X vssd1 vssd1 vccd1 vccd1 _09406_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _09335_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _09815_/A vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__buf_2
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08217_ _08217_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08372_/A sky130_fd_sc_hd__nand2_4
XFILLER_138_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09197_ _09195_/A _09195_/B _09196_/X vssd1 vssd1 vccd1 vccd1 _15574_/D sky130_fd_sc_hd__a21oi_1
XFILLER_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08148_ _07972_/A _08146_/Y _08147_/Y vssd1 vssd1 vccd1 vccd1 _08196_/A sky130_fd_sc_hd__a21o_1
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08079_ _15543_/Q vssd1 vssd1 vccd1 vccd1 _08254_/A sky130_fd_sc_hd__clkinv_2
XFILLER_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10110_ _10271_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10110_/X sky130_fd_sc_hd__or2_1
XFILLER_122_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11090_ _15924_/Q _11099_/C _10866_/X vssd1 vssd1 vccd1 vccd1 _11090_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_122_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10041_ _10082_/A _10041_/B _10041_/C vssd1 vssd1 vccd1 vccd1 _10042_/A sky130_fd_sc_hd__and3_1
XFILLER_102_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13800_ _16305_/Q _13856_/B _13800_/C vssd1 vssd1 vccd1 vccd1 _13800_/Y sky130_fd_sc_hd__nand3_1
X_11992_ _16051_/Q _12002_/C _11770_/X vssd1 vssd1 vccd1 vccd1 _11992_/Y sky130_fd_sc_hd__a21oi_1
X_14780_ _14839_/A _14780_/B _14780_/C vssd1 vssd1 vccd1 vccd1 _14781_/C sky130_fd_sc_hd__or3_1
XFILLER_44_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13731_ _16296_/Q _13731_/B _13738_/C vssd1 vssd1 vccd1 vccd1 _13733_/C sky130_fd_sc_hd__nand3_1
X_10943_ _13545_/A vssd1 vssd1 vccd1 vccd1 _11169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16450_ _16607_/CLK _16450_/D vssd1 vssd1 vccd1 vccd1 _16450_/Q sky130_fd_sc_hd__dfxtp_1
X_10874_ _15267_/B vssd1 vssd1 vccd1 vccd1 _10874_/X sky130_fd_sc_hd__buf_2
X_13662_ _13684_/C vssd1 vssd1 vccd1 vccd1 _13700_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15401_ _16101_/Q _16100_/Q _16099_/Q _15397_/X vssd1 vssd1 vccd1 vccd1 _16583_/D
+ sky130_fd_sc_hd__o31a_1
X_12613_ _16138_/Q _12776_/B _12614_/C vssd1 vssd1 vccd1 vccd1 _12613_/X sky130_fd_sc_hd__and3_1
X_16381_ _16389_/CLK _16381_/D vssd1 vssd1 vccd1 vccd1 _16381_/Q sky130_fd_sc_hd__dfxtp_1
X_13593_ _13593_/A _13600_/B vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__or2_1
X_12544_ _13392_/A vssd1 vssd1 vccd1 vccd1 _12770_/B sky130_fd_sc_hd__clkbuf_2
X_15332_ _16548_/Q _15332_/B _15335_/C vssd1 vssd1 vccd1 vccd1 _15337_/A sky130_fd_sc_hd__and3_1
X_15263_ _15260_/Y _15269_/A _15262_/Y _15258_/C vssd1 vssd1 vccd1 vccd1 _15265_/B
+ sky130_fd_sc_hd__o211a_1
X_12475_ _12495_/C vssd1 vssd1 vccd1 vccd1 _12510_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11426_ _11993_/A vssd1 vssd1 vccd1 vccd1 _11654_/B sky130_fd_sc_hd__clkbuf_2
X_14214_ _14777_/A vssd1 vssd1 vccd1 vccd1 _14439_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_6 _14113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ _16519_/Q _15247_/B _15195_/C vssd1 vssd1 vccd1 vccd1 _15194_/X sky130_fd_sc_hd__and3_1
XFILLER_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ _14145_/A _14145_/B _14145_/C vssd1 vssd1 vccd1 vccd1 _14146_/A sky130_fd_sc_hd__and3_1
X_11357_ _11357_/A vssd1 vssd1 vccd1 vccd1 _15960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10308_ _15792_/Q _10313_/B _10308_/C vssd1 vssd1 vccd1 vccd1 _10308_/Y sky130_fd_sc_hd__nand3_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14076_ _14076_/A vssd1 vssd1 vccd1 vccd1 _16344_/D sky130_fd_sc_hd__clkbuf_1
X_11288_ _11301_/C vssd1 vssd1 vccd1 vccd1 _11309_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _16197_/Q _13028_/C _12857_/X vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__a21oi_1
X_10239_ _10240_/B _10240_/C _10240_/A vssd1 vssd1 vccd1 vccd1 _10241_/B sky130_fd_sc_hd__a21o_1
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14978_ _14978_/A vssd1 vssd1 vccd1 vccd1 _16481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16717_ _16717_/A _07821_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13929_ _16325_/Q _13929_/B _13929_/C vssd1 vssd1 vccd1 vccd1 _13939_/B sky130_fd_sc_hd__and3_1
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16579_ _16595_/CLK _16579_/D vssd1 vssd1 vccd1 vccd1 _16579_/Q sky130_fd_sc_hd__dfxtp_1
X_09120_ _09076_/X _09111_/B _09115_/B _09119_/Y vssd1 vssd1 vccd1 vccd1 _15557_/D
+ sky130_fd_sc_hd__o31a_1
X_09051_ _09943_/A vssd1 vssd1 vccd1 vccd1 _09051_/X sky130_fd_sc_hd__buf_2
XFILLER_129_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08002_ _16580_/Q _08002_/B vssd1 vssd1 vccd1 vccd1 _08003_/B sky130_fd_sc_hd__or2_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09953_ _09953_/A vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__buf_2
X_08904_ _08898_/C _08899_/C _08901_/Y _08909_/A vssd1 vssd1 vccd1 vccd1 _08909_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_131_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _15713_/Q _09966_/B _09884_/C vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__and3_1
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08835_ _08835_/A _08835_/B vssd1 vssd1 vccd1 vccd1 _15495_/D sky130_fd_sc_hd__nor2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08766_ _15486_/Q _08807_/B _08766_/C vssd1 vssd1 vccd1 vccd1 _08768_/C sky130_fd_sc_hd__nand3_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08697_ _09604_/A vssd1 vssd1 vccd1 vccd1 _09117_/A sky130_fd_sc_hd__buf_2
XFILLER_53_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09318_ _09329_/C vssd1 vssd1 vccd1 vccd1 _09340_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10590_ _10590_/A vssd1 vssd1 vccd1 vccd1 _15842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09249_ _15578_/Q _15577_/Q _15576_/Q _09090_/X vssd1 vssd1 vccd1 vccd1 _15588_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ _16089_/Q _12271_/C _12036_/X vssd1 vssd1 vccd1 vccd1 _12260_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11211_ _15940_/Q _11322_/B _11211_/C vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__and3_1
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12191_ _12204_/C vssd1 vssd1 vccd1 vccd1 _12212_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11142_ _15931_/Q _11152_/C _10919_/X vssd1 vssd1 vccd1 vccd1 _11142_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15950_ _15365_/A _15950_/D vssd1 vssd1 vccd1 vccd1 _15950_/Q sky130_fd_sc_hd__dfxtp_2
X_11073_ _11088_/A _11073_/B _11073_/C vssd1 vssd1 vccd1 vccd1 _11074_/A sky130_fd_sc_hd__and3_1
XFILLER_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10024_ _15731_/Q _15730_/Q _15729_/Q _09982_/X vssd1 vssd1 vccd1 vccd1 _15741_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14901_ _16459_/Q _16458_/Q _16457_/Q _14900_/X vssd1 vssd1 vccd1 vccd1 _16469_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15881_ _16553_/Q _15881_/D vssd1 vssd1 vccd1 vccd1 _15881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14832_ _14832_/A _14839_/B vssd1 vssd1 vccd1 vccd1 _14834_/A sky130_fd_sc_hd__or2_1
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14763_ _15048_/A vssd1 vssd1 vccd1 vccd1 _14995_/B sky130_fd_sc_hd__clkbuf_2
X_11975_ _11998_/A _11975_/B _11975_/C vssd1 vssd1 vccd1 vccd1 _11976_/A sky130_fd_sc_hd__and3_1
XFILLER_72_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16502_ _16607_/CLK _16502_/D vssd1 vssd1 vccd1 vccd1 _16502_/Q sky130_fd_sc_hd__dfxtp_1
X_13714_ _13712_/A _13712_/B _13713_/X vssd1 vssd1 vccd1 vccd1 _16292_/D sky130_fd_sc_hd__a21oi_1
X_10926_ _10926_/A vssd1 vssd1 vccd1 vccd1 _15898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14694_ _14979_/A vssd1 vssd1 vccd1 vccd1 _14694_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16433_ _16595_/CLK _16433_/D vssd1 vssd1 vccd1 vccd1 _16433_/Q sky130_fd_sc_hd__dfxtp_1
X_10857_ _15891_/Q _10868_/C _10456_/A vssd1 vssd1 vccd1 vccd1 _10857_/Y sky130_fd_sc_hd__a21oi_1
X_13645_ _16285_/Q _13645_/B _13645_/C vssd1 vssd1 vccd1 vccd1 _13656_/B sky130_fd_sc_hd__and3_1
XFILLER_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _16389_/CLK _16364_/D vssd1 vssd1 vccd1 vccd1 _16364_/Q sky130_fd_sc_hd__dfxtp_1
X_10788_ _15881_/Q _10791_/C _14932_/A vssd1 vssd1 vccd1 vccd1 _10788_/Y sky130_fd_sc_hd__a21oi_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _13583_/A _13576_/B _13576_/C vssd1 vssd1 vccd1 vccd1 _13577_/A sky130_fd_sc_hd__and3_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15315_ _16710_/A _15321_/B _15315_/C vssd1 vssd1 vccd1 vccd1 _15316_/B sky130_fd_sc_hd__nand3_1
X_12527_ _12565_/A _12527_/B _12527_/C vssd1 vssd1 vccd1 vccd1 _12528_/A sky130_fd_sc_hd__and3_1
X_16295_ _16533_/Q _16295_/D vssd1 vssd1 vccd1 vccd1 _16295_/Q sky130_fd_sc_hd__dfxtp_1
X_15246_ _16528_/Q _15248_/C _10789_/B vssd1 vssd1 vccd1 vccd1 _15246_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12458_ _12455_/Y _12464_/A _12457_/Y _12453_/C vssd1 vssd1 vccd1 vccd1 _12460_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11409_ _11409_/A vssd1 vssd1 vccd1 vccd1 _15967_/D sky130_fd_sc_hd__clkbuf_1
X_15177_ _15209_/C vssd1 vssd1 vccd1 vccd1 _15215_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12389_ _12387_/Y _12383_/C _12385_/Y _12386_/X vssd1 vssd1 vccd1 vccd1 _12390_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14128_ _14126_/Y _14127_/X _14123_/C _14124_/C vssd1 vssd1 vccd1 vccd1 _14130_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14059_ _14094_/C vssd1 vssd1 vccd1 vccd1 _14101_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_141_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08620_ _08620_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _08622_/A sky130_fd_sc_hd__or2_1
X_16663__68 vssd1 vssd1 vccd1 vccd1 _16663__68/HI _16739_/A sky130_fd_sc_hd__conb_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _08548_/Y _08549_/Y _08550_/Y vssd1 vssd1 vccd1 vccd1 _15451_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08482_ _15450_/Q _08490_/A _15299_/A vssd1 vssd1 vccd1 vccd1 _08485_/A sky130_fd_sc_hd__a21o_1
XFILLER_63_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09103_ _09103_/A vssd1 vssd1 vccd1 vccd1 _15554_/D sky130_fd_sc_hd__clkbuf_1
X_09034_ _09029_/B _09032_/B _08914_/X vssd1 vssd1 vccd1 vccd1 _09042_/C sky130_fd_sc_hd__o21a_1
XFILLER_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09936_ _08654_/X _09932_/B _09792_/X vssd1 vssd1 vccd1 vccd1 _09938_/A sky130_fd_sc_hd__a21oi_1
XFILLER_132_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09867_ _15710_/Q _09867_/B _09873_/C vssd1 vssd1 vccd1 vccd1 _09869_/C sky130_fd_sc_hd__nand3_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08818_ input3/X vssd1 vssd1 vccd1 vccd1 _14806_/A sky130_fd_sc_hd__buf_4
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09798_ _09816_/C vssd1 vssd1 vccd1 vccd1 _09836_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _09294_/A vssd1 vssd1 vccd1 vccd1 _08921_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11760_ _11776_/A _11760_/B _11760_/C vssd1 vssd1 vccd1 vccd1 _11761_/A sky130_fd_sc_hd__and3_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10759_/A _10711_/B vssd1 vssd1 vccd1 vccd1 _10711_/X sky130_fd_sc_hd__or2_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11691_ _16008_/Q _11750_/B _11698_/C vssd1 vssd1 vccd1 vccd1 _11693_/C sky130_fd_sc_hd__nand3_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _10649_/A _10642_/B _10642_/C vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__and3_1
X_13430_ _13598_/A vssd1 vssd1 vccd1 vccd1 _13470_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _13359_/Y _13354_/C _13356_/Y _13366_/A vssd1 vssd1 vccd1 vccd1 _13366_/B
+ sky130_fd_sc_hd__a211oi_1
X_10573_ _10573_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _10573_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15100_ _15100_/A _15100_/B _15100_/C vssd1 vssd1 vccd1 vccd1 _15101_/A sky130_fd_sc_hd__and3_1
X_12312_ _12312_/A vssd1 vssd1 vccd1 vccd1 _12535_/B sky130_fd_sc_hd__clkbuf_2
X_16080_ _16118_/CLK _16080_/D vssd1 vssd1 vccd1 vccd1 _16080_/Q sky130_fd_sc_hd__dfxtp_1
X_13292_ _16233_/Q _13292_/B _13292_/C vssd1 vssd1 vccd1 vccd1 _13292_/Y sky130_fd_sc_hd__nand3_1
X_12243_ _12304_/A _12243_/B _12243_/C vssd1 vssd1 vccd1 vccd1 _12244_/C sky130_fd_sc_hd__or3_1
X_15031_ _15031_/A vssd1 vssd1 vccd1 vccd1 _16490_/D sky130_fd_sc_hd__clkbuf_1
X_12174_ _16075_/Q _12347_/B _12179_/C vssd1 vssd1 vccd1 vccd1 _12174_/Y sky130_fd_sc_hd__nand3_1
X_11125_ _11125_/A vssd1 vssd1 vccd1 vccd1 _15927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15933_ _15365_/A _15933_/D vssd1 vssd1 vccd1 vccd1 _15933_/Q sky130_fd_sc_hd__dfxtp_1
X_11056_ _16561_/Q vssd1 vssd1 vccd1 vccd1 _11070_/C sky130_fd_sc_hd__inv_2
X_10007_ _10005_/A _10005_/B _10004_/Y _10006_/Y vssd1 vssd1 vccd1 vccd1 _15736_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15864_ _16570_/CLK _15864_/D vssd1 vssd1 vccd1 vccd1 _15864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14815_ _16457_/Q _15041_/B _14823_/C vssd1 vssd1 vccd1 vccd1 _14815_/X sky130_fd_sc_hd__and3_1
X_15795_ _16595_/CLK _15795_/D vssd1 vssd1 vccd1 vccd1 _15795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14746_ _14746_/A vssd1 vssd1 vccd1 vccd1 _16445_/D sky130_fd_sc_hd__clkbuf_1
X_11958_ _12185_/A vssd1 vssd1 vccd1 vccd1 _11998_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10909_ _10902_/C _10903_/C _10906_/Y _10907_/X vssd1 vssd1 vccd1 vccd1 _10910_/C
+ sky130_fd_sc_hd__a211o_1
X_14677_ _14697_/C vssd1 vssd1 vccd1 vccd1 _14710_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11889_ _11889_/A vssd1 vssd1 vccd1 vccd1 _16034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16416_ input11/X _16416_/D vssd1 vssd1 vccd1 vccd1 _16416_/Q sky130_fd_sc_hd__dfxtp_2
X_13628_ _13635_/A _13628_/B _13628_/C vssd1 vssd1 vccd1 vccd1 _13629_/A sky130_fd_sc_hd__and3_1
XFILLER_13_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16347_ _16389_/CLK _16347_/D vssd1 vssd1 vccd1 vccd1 _16347_/Q sky130_fd_sc_hd__dfxtp_1
X_13559_ _16272_/Q _13731_/B _13565_/C vssd1 vssd1 vccd1 vccd1 _13561_/C sky130_fd_sc_hd__nand3_1
XFILLER_146_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16278_ _16533_/Q _16278_/D vssd1 vssd1 vccd1 vccd1 _16278_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15229_ _15248_/C vssd1 vssd1 vccd1 vccd1 _15261_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07982_ _07982_/A _07982_/B vssd1 vssd1 vccd1 vccd1 _07983_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09721_ _09722_/B _09722_/C _09722_/A vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__a21o_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09652_ _09647_/Y _09650_/X _09651_/X vssd1 vssd1 vccd1 vccd1 _09652_/Y sky130_fd_sc_hd__a21oi_1
X_08603_ _10294_/C vssd1 vssd1 vccd1 vccd1 _08604_/A sky130_fd_sc_hd__clkbuf_2
X_09583_ _10183_/A vssd1 vssd1 vccd1 vccd1 _09583_/X sky130_fd_sc_hd__buf_2
XFILLER_103_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ _08516_/B _08534_/B vssd1 vssd1 vccd1 vccd1 _08556_/A sky130_fd_sc_hd__and2b_1
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08465_ _08466_/A _08466_/B vssd1 vssd1 vccd1 vccd1 _08502_/A sky130_fd_sc_hd__or2_1
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08396_ _08396_/A _08396_/B vssd1 vssd1 vccd1 vccd1 _08396_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09017_ _09018_/B _09018_/C _09018_/A vssd1 vssd1 vccd1 vccd1 _09019_/B sky130_fd_sc_hd__a21o_1
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09919_ _15721_/Q _09919_/B _09925_/C vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__and3_1
X_12930_ _12952_/C vssd1 vssd1 vccd1 vccd1 _12967_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12861_/A _12868_/B vssd1 vssd1 vccd1 vccd1 _12863_/A sky130_fd_sc_hd__or2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14598_/Y _14594_/C _14596_/Y _14605_/A vssd1 vssd1 vccd1 vccd1 _14605_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11812_/A vssd1 vssd1 vccd1 vccd1 _16023_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _16551_/CLK _15580_/D vssd1 vssd1 vccd1 vccd1 _15580_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _16164_/Q _13022_/B _12792_/C vssd1 vssd1 vccd1 vccd1 _12800_/A sky130_fd_sc_hd__and3_1
XFILLER_26_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _16412_/Q _14756_/B _14539_/C vssd1 vssd1 vccd1 vccd1 _14531_/X sky130_fd_sc_hd__and3_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11779_/C vssd1 vssd1 vccd1 vccd1 _11785_/C sky130_fd_sc_hd__clkbuf_2
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14462_ _14462_/A vssd1 vssd1 vccd1 vccd1 _16400_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11901_/A _11679_/C vssd1 vssd1 vccd1 vccd1 _11674_/X sky130_fd_sc_hd__or2_1
X_16201_ _16555_/Q _16201_/D vssd1 vssd1 vccd1 vccd1 _16201_/Q sky130_fd_sc_hd__dfxtp_1
X_13413_ _13413_/A vssd1 vssd1 vccd1 vccd1 _16250_/D sky130_fd_sc_hd__clkbuf_1
X_10625_ _15867_/Q vssd1 vssd1 vccd1 vccd1 _10630_/C sky130_fd_sc_hd__inv_2
X_14393_ _14406_/C vssd1 vssd1 vccd1 vccd1 _14414_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16132_ _16554_/Q _16132_/D vssd1 vssd1 vccd1 vccd1 _16132_/Q sky130_fd_sc_hd__dfxtp_1
X_10556_ _10589_/A _10556_/B _10556_/C vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__and3_1
X_13344_ _16241_/Q _13573_/B _13344_/C vssd1 vssd1 vccd1 vccd1 _13344_/Y sky130_fd_sc_hd__nand3_1
XFILLER_10_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16063_ _16118_/CLK _16063_/D vssd1 vssd1 vccd1 vccd1 _16063_/Q sky130_fd_sc_hd__dfxtp_1
X_13275_ _13362_/A _13275_/B _13279_/A vssd1 vssd1 vccd1 vccd1 _16230_/D sky130_fd_sc_hd__nor3_1
X_10487_ _15826_/Q _10679_/B _10494_/C vssd1 vssd1 vccd1 vccd1 _10489_/C sky130_fd_sc_hd__nand3_1
XFILLER_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15014_ _15027_/C vssd1 vssd1 vccd1 vccd1 _15035_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12226_ _16084_/Q _12456_/B _12226_/C vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__and3_1
XFILLER_69_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12157_ _13006_/A vssd1 vssd1 vccd1 vccd1 _12157_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _11109_/B _11109_/C _10999_/X vssd1 vssd1 vccd1 vccd1 _11110_/B sky130_fd_sc_hd__o21ai_1
XFILLER_150_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12088_ _12089_/B _12089_/C _12089_/A vssd1 vssd1 vccd1 vccd1 _12090_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15916_ _15365_/A _15916_/D vssd1 vssd1 vccd1 vccd1 _15916_/Q sky130_fd_sc_hd__dfxtp_1
X_11039_ _15916_/Q _11039_/B _11039_/C vssd1 vssd1 vccd1 vccd1 _11047_/A sky130_fd_sc_hd__and3_1
XFILLER_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16633__38 vssd1 vssd1 vccd1 vccd1 _16633__38/HI _16699_/A sky130_fd_sc_hd__conb_1
XFILLER_94_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15847_ _16551_/CLK _15847_/D vssd1 vssd1 vccd1 vccd1 _15847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15778_ _16595_/CLK _15778_/D vssd1 vssd1 vccd1 vccd1 _15778_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14729_ _14742_/C vssd1 vssd1 vccd1 vccd1 _14750_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_08250_ _08251_/A _08251_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08252_/A sky130_fd_sc_hd__a21oi_1
XFILLER_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08181_ _08181_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08181_/X sky130_fd_sc_hd__or2_1
XFILLER_146_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07965_ _13777_/A _07965_/B vssd1 vssd1 vccd1 vccd1 _08181_/B sky130_fd_sc_hd__xnor2_2
XFILLER_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09704_ _09529_/X _09701_/B _09703_/Y vssd1 vssd1 vccd1 vccd1 _15676_/D sky130_fd_sc_hd__o21a_1
XFILLER_68_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07896_ _09255_/C _07896_/B vssd1 vssd1 vccd1 vccd1 _08116_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09635_ _15666_/Q _09636_/C _09590_/X vssd1 vssd1 vccd1 vccd1 _09635_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09566_ _09560_/Y _09561_/X _09563_/B vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__o21a_1
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08517_ _08532_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__xor2_2
X_09497_ _09497_/A _09497_/B _09501_/A vssd1 vssd1 vccd1 vccd1 _15634_/D sky130_fd_sc_hd__nor3_1
XFILLER_70_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08448_ _08379_/B _08448_/B vssd1 vssd1 vccd1 vccd1 _08449_/B sky130_fd_sc_hd__and2b_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _08448_/B _08379_/B vssd1 vssd1 vccd1 vccd1 _08399_/A sky130_fd_sc_hd__xnor2_4
XFILLER_137_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10410_ _10410_/A _10410_/B vssd1 vssd1 vccd1 vccd1 _10411_/B sky130_fd_sc_hd__nor2_1
X_11390_ _11391_/B _11391_/C _11282_/X vssd1 vssd1 vccd1 vccd1 _11392_/B sky130_fd_sc_hd__o21ai_1
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ _15800_/Q _10342_/C _10243_/X vssd1 vssd1 vccd1 vccd1 _10341_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ _13060_/A vssd1 vssd1 vccd1 vccd1 _14186_/A sky130_fd_sc_hd__buf_4
X_10272_ _10270_/A _10270_/B _10271_/X vssd1 vssd1 vccd1 vccd1 _15783_/D sky130_fd_sc_hd__a21oi_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12011_ _12011_/A _12018_/B vssd1 vssd1 vccd1 vccd1 _12013_/A sky130_fd_sc_hd__or2_1
XFILLER_3_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16750_ _16750_/A _07767_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
X_13962_ _13962_/A vssd1 vssd1 vccd1 vccd1 _16328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _15791_/CLK _15701_/D vssd1 vssd1 vccd1 vccd1 _15701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12913_ _12911_/Y _12907_/C _12909_/Y _12918_/A vssd1 vssd1 vccd1 vccd1 _12918_/B
+ sky130_fd_sc_hd__a211oi_1
X_13893_ _16320_/Q _13900_/C _13729_/X vssd1 vssd1 vccd1 vccd1 _13896_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15632_ _15812_/CLK _15632_/D vssd1 vssd1 vccd1 vccd1 _15632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12844_ _16170_/Q _12904_/B _12852_/C vssd1 vssd1 vccd1 vccd1 _12844_/Y sky130_fd_sc_hd__nand3_1
XFILLER_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15791_/CLK _15563_/D vssd1 vssd1 vccd1 vccd1 _15563_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _16162_/Q _12778_/C _12723_/X vssd1 vssd1 vccd1 vccd1 _12775_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _16410_/Q _14524_/C _14294_/X vssd1 vssd1 vccd1 vccd1 _14514_/Y sky130_fd_sc_hd__a21oi_1
X_11726_ _12292_/A vssd1 vssd1 vccd1 vccd1 _11726_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _16570_/CLK _15494_/D vssd1 vssd1 vccd1 vccd1 _15494_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14445_ _14458_/C vssd1 vssd1 vccd1 vccd1 _14466_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11657_ _11655_/Y _11651_/C _11653_/Y _11654_/X vssd1 vssd1 vccd1 vccd1 _11658_/C
+ sky130_fd_sc_hd__a211o_1
X_10608_ _10605_/Y _10614_/A _10607_/Y _10603_/C vssd1 vssd1 vccd1 vccd1 _10610_/B
+ sky130_fd_sc_hd__o211a_1
X_14376_ _14372_/Y _14382_/A _14375_/Y _14369_/C vssd1 vssd1 vccd1 vccd1 _14378_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11588_ _11582_/C _11583_/C _11585_/Y _11586_/X vssd1 vssd1 vccd1 vccd1 _11589_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_143_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16115_ _16554_/Q _16115_/D vssd1 vssd1 vccd1 vccd1 _16115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13327_ _16239_/Q _13383_/B _13336_/C vssd1 vssd1 vccd1 vccd1 _13332_/A sky130_fd_sc_hd__and3_1
XFILLER_143_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10539_ _15835_/Q _10679_/B _10546_/C vssd1 vssd1 vccd1 vccd1 _10541_/C sky130_fd_sc_hd__nand3_1
XFILLER_142_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _16118_/CLK _16046_/D vssd1 vssd1 vccd1 vccd1 _16046_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13258_ _13258_/A _13266_/B vssd1 vssd1 vccd1 vccd1 _13260_/A sky130_fd_sc_hd__or2_1
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12209_ _16082_/Q _12212_/C _12157_/X vssd1 vssd1 vccd1 vccd1 _12209_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13189_ _13187_/Y _13181_/C _13185_/Y _13186_/X vssd1 vssd1 vccd1 vccd1 _13190_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09420_ _15622_/Q _09428_/C _10750_/B vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__a21oi_1
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ _10418_/A vssd1 vssd1 vccd1 vccd1 _09351_/X sky130_fd_sc_hd__clkbuf_2
X_08302_ _08302_/A vssd1 vssd1 vccd1 vccd1 _08849_/C sky130_fd_sc_hd__clkbuf_2
X_09282_ _09277_/A _09276_/Y _09277_/B vssd1 vssd1 vccd1 vccd1 _09282_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_33_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08233_ _10332_/C _08035_/B _08034_/A vssd1 vssd1 vccd1 vccd1 _08380_/A sky130_fd_sc_hd__o21ai_4
XFILLER_119_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08164_ _08165_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__nor2_1
XFILLER_118_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08095_ _15696_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08096_/B sky130_fd_sc_hd__xnor2_1
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08997_ _08992_/B _08995_/B _08914_/X vssd1 vssd1 vccd1 vccd1 _09003_/C sky130_fd_sc_hd__o21a_1
XFILLER_88_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07948_ _07948_/A _07948_/B vssd1 vssd1 vccd1 vccd1 _07949_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07879_ _16424_/Q _16406_/Q vssd1 vssd1 vccd1 vccd1 _08129_/A sky130_fd_sc_hd__nand2_2
XFILLER_28_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09618_ _09617_/X _09486_/X _09611_/B _09487_/X vssd1 vssd1 vccd1 vccd1 _09619_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _10907_/C vssd1 vssd1 vccd1 vccd1 _10914_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09549_ _15648_/Q _09550_/C _09369_/X vssd1 vssd1 vccd1 vccd1 _09549_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12560_ _13407_/A vssd1 vssd1 vccd1 vccd1 _12784_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _11511_/A vssd1 vssd1 vccd1 vccd1 _15981_/D sky130_fd_sc_hd__clkbuf_1
X_12491_ _12491_/A vssd1 vssd1 vccd1 vccd1 _16120_/D sky130_fd_sc_hd__clkbuf_1
X_14230_ _16368_/Q _14289_/B _14237_/C vssd1 vssd1 vccd1 vccd1 _14232_/C sky130_fd_sc_hd__nand3_1
X_11442_ _15973_/Q _11444_/C _11441_/X vssd1 vssd1 vccd1 vccd1 _11445_/A sky130_fd_sc_hd__a21oi_1
XFILLER_109_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ _15964_/Q _11381_/C _11150_/X vssd1 vssd1 vccd1 vccd1 _11373_/Y sky130_fd_sc_hd__a21oi_1
X_14161_ _14162_/B _14162_/C _14108_/X vssd1 vssd1 vccd1 vccd1 _14163_/B sky130_fd_sc_hd__o21ai_1
X_10324_ _10168_/X _10322_/B _10224_/X vssd1 vssd1 vccd1 vccd1 _10324_/Y sky130_fd_sc_hd__a21oi_1
X_13112_ _16209_/Q _13336_/B _13112_/C vssd1 vssd1 vccd1 vccd1 _13112_/X sky130_fd_sc_hd__and3_1
X_14092_ _14092_/A vssd1 vssd1 vccd1 vccd1 _14205_/A sky130_fd_sc_hd__buf_2
XFILLER_124_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10255_ _15782_/Q _10396_/B _10261_/C vssd1 vssd1 vccd1 vccd1 _10255_/Y sky130_fd_sc_hd__nand3_1
X_13043_ _16199_/Q _13082_/C _12933_/X vssd1 vssd1 vccd1 vccd1 _13045_/B sky130_fd_sc_hd__a21oi_1
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10186_ _10186_/A _10186_/B _10186_/C vssd1 vssd1 vccd1 vccd1 _10187_/C sky130_fd_sc_hd__nand3_1
XFILLER_94_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14994_ _16485_/Q _15001_/C _14821_/X vssd1 vssd1 vccd1 vccd1 _14994_/Y sky130_fd_sc_hd__a21oi_1
X_16733_ _16733_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _13966_/C vssd1 vssd1 vccd1 vccd1 _13981_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13876_ _13876_/A _13883_/B vssd1 vssd1 vccd1 vccd1 _13878_/A sky130_fd_sc_hd__or2_1
XFILLER_35_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15615_ _16570_/CLK _15615_/D vssd1 vssd1 vccd1 vccd1 _15615_/Q sky130_fd_sc_hd__dfxtp_1
X_12827_ _13392_/A vssd1 vssd1 vccd1 vccd1 _13053_/B sky130_fd_sc_hd__clkbuf_2
X_16595_ _16595_/CLK _16595_/D vssd1 vssd1 vccd1 vccd1 _16595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15546_ _15791_/CLK _15546_/D vssd1 vssd1 vccd1 vccd1 _15546_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12778_/C vssd1 vssd1 vccd1 vccd1 _12792_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _11717_/A _11709_/B _11709_/C vssd1 vssd1 vccd1 vccd1 _11710_/A sky130_fd_sc_hd__and3_1
X_15477_ _16570_/CLK _15477_/D vssd1 vssd1 vccd1 vccd1 _15477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12689_ _12687_/Y _12681_/C _12684_/Y _12694_/A vssd1 vssd1 vccd1 vccd1 _12694_/B
+ sky130_fd_sc_hd__a211oi_1
X_14428_ _16395_/Q _14598_/B _14433_/C vssd1 vssd1 vccd1 vccd1 _14428_/Y sky130_fd_sc_hd__nand3_1
XFILLER_128_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14359_ _14356_/Y _14357_/X _14358_/Y _14354_/C vssd1 vssd1 vccd1 vccd1 _14361_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08920_ _08920_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _15513_/D sky130_fd_sc_hd__nor2_1
X_16029_ _16554_/Q _16029_/D vssd1 vssd1 vccd1 vccd1 _16029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08851_ _08851_/A _08851_/B _08851_/C vssd1 vssd1 vccd1 vccd1 _08852_/C sky130_fd_sc_hd__nand3_1
XFILLER_112_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07802_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07802_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08782_ _08782_/A _08782_/B vssd1 vssd1 vccd1 vccd1 _08783_/B sky130_fd_sc_hd__nor2_1
XFILLER_111_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09403_ _09416_/C vssd1 vssd1 vccd1 vccd1 _09428_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09334_ _15604_/Q _09837_/A _09340_/C vssd1 vssd1 vccd1 vccd1 _09336_/B sky130_fd_sc_hd__and3_1
XFILLER_139_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09265_ _15594_/Q _09267_/C _15341_/B vssd1 vssd1 vccd1 vccd1 _09265_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08216_ _14444_/A _08036_/B _08039_/A vssd1 vssd1 vccd1 vccd1 _08220_/A sky130_fd_sc_hd__o21ai_4
X_09196_ _09849_/A _09196_/B vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__or2_1
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08147_ _09802_/C _08147_/B vssd1 vssd1 vccd1 vccd1 _08147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08078_ _14902_/A _08248_/B vssd1 vssd1 vccd1 vccd1 _08090_/A sky130_fd_sc_hd__xnor2_4
XFILLER_134_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16669__74 vssd1 vssd1 vccd1 vccd1 _16669__74/HI _16745_/A sky130_fd_sc_hd__conb_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _10034_/C _10035_/C _10037_/Y _10038_/X vssd1 vssd1 vccd1 vccd1 _10041_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11991_ _11991_/A vssd1 vssd1 vccd1 vccd1 _16049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _16296_/Q _13738_/C _13729_/X vssd1 vssd1 vccd1 vccd1 _13733_/B sky130_fd_sc_hd__a21o_1
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10942_ input7/X vssd1 vssd1 vccd1 vccd1 _13545_/A sky130_fd_sc_hd__buf_6
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ _13676_/C vssd1 vssd1 vccd1 vccd1 _13684_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10873_ _12574_/A vssd1 vssd1 vccd1 vccd1 _15267_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15400_ _16093_/Q _16092_/Q _16091_/Q _15397_/X vssd1 vssd1 vccd1 vccd1 _16582_/D
+ sky130_fd_sc_hd__o31a_1
X_12612_ _16138_/Q _12614_/C _12440_/X vssd1 vssd1 vccd1 vccd1 _12612_/Y sky130_fd_sc_hd__a21oi_1
X_16380_ _16389_/CLK _16380_/D vssd1 vssd1 vccd1 vccd1 _16380_/Q sky130_fd_sc_hd__dfxtp_1
X_13592_ _16277_/Q _13645_/B _13592_/C vssd1 vssd1 vccd1 vccd1 _13600_/B sky130_fd_sc_hd__and3_1
X_15331_ _16548_/Q _15346_/C _08843_/A vssd1 vssd1 vccd1 vccd1 _15333_/B sky130_fd_sc_hd__a21oi_1
XFILLER_40_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12543_ _16129_/Q _12554_/C _12323_/X vssd1 vssd1 vccd1 vccd1 _12543_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15262_ _16529_/Q _15262_/B _15267_/C vssd1 vssd1 vccd1 vccd1 _15262_/Y sky130_fd_sc_hd__nand3_1
X_12474_ _12487_/C vssd1 vssd1 vccd1 vccd1 _12495_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14213_ _14211_/A _14211_/B _14212_/X vssd1 vssd1 vccd1 vccd1 _16364_/D sky130_fd_sc_hd__a21oi_1
X_11425_ _15971_/Q _11436_/C _11202_/X vssd1 vssd1 vccd1 vccd1 _11425_/Y sky130_fd_sc_hd__a21oi_1
X_15193_ _16519_/Q _15195_/C _14979_/X vssd1 vssd1 vccd1 vccd1 _15193_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_7 _14113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14144_ _14142_/Y _14138_/C _14140_/Y _14141_/X vssd1 vssd1 vccd1 vccd1 _14145_/C
+ sky130_fd_sc_hd__a211o_1
X_11356_ _11371_/A _11356_/B _11356_/C vssd1 vssd1 vccd1 vccd1 _11357_/A sky130_fd_sc_hd__and3_1
XFILLER_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ _15793_/Q _10307_/B _10307_/C vssd1 vssd1 vccd1 vccd1 _10315_/A sky130_fd_sc_hd__and3_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14075_ _14090_/A _14075_/B _14075_/C vssd1 vssd1 vccd1 vccd1 _14076_/A sky130_fd_sc_hd__and3_1
X_11287_ _11287_/A vssd1 vssd1 vccd1 vccd1 _11301_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _13080_/A _13026_/B _13030_/B vssd1 vssd1 vccd1 vccd1 _16195_/D sky130_fd_sc_hd__nor3_1
X_10238_ _15781_/Q _10434_/B _10247_/C vssd1 vssd1 vccd1 vccd1 _10240_/C sky130_fd_sc_hd__nand3_1
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10169_ _10168_/X _10166_/B _10012_/X vssd1 vssd1 vccd1 vccd1 _10169_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14977_ _14992_/A _14977_/B _14977_/C vssd1 vssd1 vccd1 vccd1 _14978_/A sky130_fd_sc_hd__and3_1
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16716_ _16716_/A _07820_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_81_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13928_ _16325_/Q _13929_/C _13705_/X vssd1 vssd1 vccd1 vccd1 _13930_/A sky130_fd_sc_hd__a21oi_1
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13859_ _13866_/A _13859_/B _13859_/C vssd1 vssd1 vccd1 vccd1 _13860_/A sky130_fd_sc_hd__and3_1
XFILLER_23_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16578_ _16595_/CLK _16578_/D vssd1 vssd1 vccd1 vccd1 _16578_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_148_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15529_ _15791_/CLK _15529_/D vssd1 vssd1 vccd1 vccd1 _15529_/Q sky130_fd_sc_hd__dfxtp_2
X_09050_ _14906_/A vssd1 vssd1 vccd1 vccd1 _09943_/A sky130_fd_sc_hd__clkbuf_4
X_08001_ _16580_/Q _08002_/B vssd1 vssd1 vccd1 vccd1 _08003_/A sky130_fd_sc_hd__nand2_1
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09952_ _09952_/A vssd1 vssd1 vccd1 vccd1 _15725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08903_ _08901_/Y _08909_/A _08898_/C _08899_/C vssd1 vssd1 vccd1 vccd1 _08905_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09880_/A _09879_/Y _09880_/B vssd1 vssd1 vccd1 vccd1 _09883_/Y sky130_fd_sc_hd__o21bai_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08832_/X _08836_/C _08833_/X vssd1 vssd1 vccd1 vccd1 _08835_/B sky130_fd_sc_hd__o21ai_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _15486_/Q _08766_/C _15335_/B vssd1 vssd1 vccd1 vccd1 _08768_/B sky130_fd_sc_hd__a21o_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08696_ _10456_/A vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09317_ _09320_/C vssd1 vssd1 vccd1 vccd1 _09329_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_09248_ _09087_/X _09246_/A _09247_/Y vssd1 vssd1 vccd1 vccd1 _15587_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09179_ _09180_/B _09180_/C _09180_/A vssd1 vssd1 vccd1 vccd1 _09181_/B sky130_fd_sc_hd__a21o_1
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11210_ _15940_/Q _11217_/C _11150_/X vssd1 vssd1 vccd1 vccd1 _11210_/Y sky130_fd_sc_hd__a21oi_1
X_12190_ _16581_/Q vssd1 vssd1 vccd1 vccd1 _12204_/C sky130_fd_sc_hd__inv_2
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11141_ _11141_/A vssd1 vssd1 vccd1 vccd1 _15929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11072_ _11066_/C _11067_/C _11069_/Y _11070_/X vssd1 vssd1 vccd1 vccd1 _11073_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10023_ _10023_/A _10023_/B vssd1 vssd1 vccd1 vccd1 _15740_/D sky130_fd_sc_hd__nor2_1
X_14900_ _15378_/A vssd1 vssd1 vccd1 vccd1 _14900_/X sky130_fd_sc_hd__buf_2
XFILLER_49_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15880_ _16553_/Q _15880_/D vssd1 vssd1 vccd1 vccd1 _15880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14831_ _16459_/Q _15055_/B _14831_/C vssd1 vssd1 vccd1 vccd1 _14839_/B sky130_fd_sc_hd__and3_1
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14762_ _16449_/Q _14770_/C _14537_/X vssd1 vssd1 vccd1 vccd1 _14762_/Y sky130_fd_sc_hd__a21oi_1
X_11974_ _11974_/A _11974_/B _11974_/C vssd1 vssd1 vccd1 vccd1 _11975_/C sky130_fd_sc_hd__nand3_1
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16501_ _16607_/CLK _16501_/D vssd1 vssd1 vccd1 vccd1 _16501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13713_ _13879_/A _13717_/C vssd1 vssd1 vccd1 vccd1 _13713_/X sky130_fd_sc_hd__or2_1
X_10925_ _10925_/A _10925_/B _10925_/C vssd1 vssd1 vccd1 vccd1 _10926_/A sky130_fd_sc_hd__and3_1
XFILLER_17_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14693_ _14693_/A vssd1 vssd1 vccd1 vccd1 _16436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16432_ _16607_/CLK _16432_/D vssd1 vssd1 vccd1 vccd1 _16432_/Q sky130_fd_sc_hd__dfxtp_1
X_13644_ _16285_/Q _13645_/C _13421_/X vssd1 vssd1 vccd1 vccd1 _13646_/A sky130_fd_sc_hd__a21oi_1
X_10856_ _10856_/A vssd1 vssd1 vccd1 vccd1 _15889_/D sky130_fd_sc_hd__clkbuf_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16389_/CLK _16363_/D vssd1 vssd1 vccd1 vccd1 _16363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13573_/Y _13568_/C _13571_/Y _13572_/X vssd1 vssd1 vccd1 vccd1 _13576_/C
+ sky130_fd_sc_hd__a211o_1
X_10787_ _14979_/A vssd1 vssd1 vccd1 vccd1 _14932_/A sky130_fd_sc_hd__clkbuf_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _16710_/A _15321_/B _15315_/C vssd1 vssd1 vccd1 vccd1 _15320_/A sky130_fd_sc_hd__a21o_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _12586_/A _12526_/B _12526_/C vssd1 vssd1 vccd1 vccd1 _12527_/C sky130_fd_sc_hd__or3_1
X_16294_ _16533_/Q _16294_/D vssd1 vssd1 vccd1 vccd1 _16294_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15245_ _15245_/A vssd1 vssd1 vccd1 vccd1 _16526_/D sky130_fd_sc_hd__clkbuf_1
X_12457_ _16115_/Q _12629_/B _12462_/C vssd1 vssd1 vccd1 vccd1 _12457_/Y sky130_fd_sc_hd__nand3_1
X_11408_ _11431_/A _11408_/B _11408_/C vssd1 vssd1 vccd1 vccd1 _11409_/A sky130_fd_sc_hd__and3_1
X_15176_ _15195_/C vssd1 vssd1 vccd1 vccd1 _15209_/C sky130_fd_sc_hd__clkbuf_1
X_12388_ _12385_/Y _12386_/X _12387_/Y _12383_/C vssd1 vssd1 vccd1 vccd1 _12390_/B
+ sky130_fd_sc_hd__o211ai_1
X_14127_ _16353_/Q _14179_/B _14127_/C vssd1 vssd1 vccd1 vccd1 _14127_/X sky130_fd_sc_hd__and3_1
X_11339_ _11339_/A vssd1 vssd1 vccd1 vccd1 _11353_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14058_ _14079_/C vssd1 vssd1 vccd1 vccd1 _14094_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13009_ _16193_/Q _13009_/B _13009_/C vssd1 vssd1 vccd1 vccd1 _13009_/Y sky130_fd_sc_hd__nand3_1
XFILLER_121_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08550_ _08548_/Y _08549_/Y _15344_/A vssd1 vssd1 vccd1 vccd1 _08550_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08481_ _08481_/A _08481_/B vssd1 vssd1 vccd1 vccd1 _15299_/A sky130_fd_sc_hd__xnor2_2
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09102_ _09142_/A _09102_/B _09102_/C vssd1 vssd1 vccd1 vccd1 _09103_/A sky130_fd_sc_hd__and3_1
XFILLER_148_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09033_ _09031_/A _09031_/B _09032_/X vssd1 vssd1 vccd1 vccd1 _15538_/D sky130_fd_sc_hd__a21oi_1
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09935_ _09749_/X _09932_/B _09934_/Y vssd1 vssd1 vccd1 vccd1 _15721_/D sky130_fd_sc_hd__o21a_1
X_16639__44 vssd1 vssd1 vccd1 vccd1 _16639__44/HI _16715_/A sky130_fd_sc_hd__conb_1
XFILLER_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _15710_/Q _09873_/C _08589_/A vssd1 vssd1 vccd1 vccd1 _09869_/B sky130_fd_sc_hd__a21o_1
XFILLER_100_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _15497_/Q _08822_/C _08777_/X vssd1 vssd1 vccd1 vccd1 _08823_/A sky130_fd_sc_hd__a21oi_1
X_09797_ _09802_/C vssd1 vssd1 vccd1 vccd1 _09816_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _08748_/A vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _08680_/B _08680_/C _08680_/A vssd1 vssd1 vccd1 vccd1 _08681_/B sky130_fd_sc_hd__a21o_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10710_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10711_/B sky130_fd_sc_hd__nor2_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _16008_/Q _11698_/C _11463_/X vssd1 vssd1 vccd1 vccd1 _11693_/B sky130_fd_sc_hd__a21o_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ _10635_/C _10636_/C _10638_/Y _10639_/X vssd1 vssd1 vccd1 vccd1 _10642_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13360_ _13356_/Y _13366_/A _13359_/Y _13354_/C vssd1 vssd1 vccd1 vccd1 _13362_/B
+ sky130_fd_sc_hd__o211a_1
X_10572_ _10566_/B _10570_/B _10414_/X vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__o21a_1
X_12311_ _16095_/Q _12352_/C _12081_/X vssd1 vssd1 vccd1 vccd1 _12314_/B sky130_fd_sc_hd__a21oi_1
XFILLER_139_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13291_ _16234_/Q _13342_/B _13292_/C vssd1 vssd1 vccd1 vccd1 _13291_/X sky130_fd_sc_hd__and3_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15030_ _15045_/A _15030_/B _15030_/C vssd1 vssd1 vccd1 vccd1 _15031_/A sky130_fd_sc_hd__and3_1
XFILLER_142_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12242_ _12243_/B _12243_/C _12133_/X vssd1 vssd1 vccd1 vccd1 _12244_/B sky130_fd_sc_hd__o21ai_1
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _16076_/Q _12173_/B _12173_/C vssd1 vssd1 vccd1 vccd1 _12181_/A sky130_fd_sc_hd__and3_1
X_11124_ _11148_/A _11124_/B _11124_/C vssd1 vssd1 vccd1 vccd1 _11125_/A sky130_fd_sc_hd__and3_1
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15932_ _15365_/A _15932_/D vssd1 vssd1 vccd1 vccd1 _15932_/Q sky130_fd_sc_hd__dfxtp_1
X_11055_ _11055_/A vssd1 vssd1 vccd1 vccd1 _15917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _10005_/X _10004_/Y _08700_/A vssd1 vssd1 vccd1 vccd1 _10006_/Y sky130_fd_sc_hd__a21oi_1
X_15863_ _16570_/CLK _15863_/D vssd1 vssd1 vccd1 vccd1 _15863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14814_ _14814_/A vssd1 vssd1 vccd1 vccd1 _15041_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_91_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15794_ _15812_/CLK _15794_/D vssd1 vssd1 vccd1 vccd1 _15794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14745_ _14760_/A _14745_/B _14745_/C vssd1 vssd1 vccd1 vccd1 _14746_/A sky130_fd_sc_hd__and3_1
X_11957_ _11957_/A vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ _10906_/Y _10907_/X _10902_/C _10903_/C vssd1 vssd1 vccd1 vccd1 _10910_/B
+ sky130_fd_sc_hd__o211ai_1
X_14676_ _14689_/C vssd1 vssd1 vccd1 vccd1 _14697_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11888_ _11888_/A _11888_/B _11888_/C vssd1 vssd1 vccd1 vccd1 _11889_/A sky130_fd_sc_hd__and3_1
X_16415_ input11/X _16415_/D vssd1 vssd1 vccd1 vccd1 _16415_/Q sky130_fd_sc_hd__dfxtp_1
X_13627_ _13625_/Y _13620_/C _13622_/Y _13623_/X vssd1 vssd1 vccd1 vccd1 _13628_/C
+ sky130_fd_sc_hd__a211o_1
X_10839_ _10864_/A _10839_/B _10839_/C vssd1 vssd1 vccd1 vccd1 _10840_/A sky130_fd_sc_hd__and3_1
XFILLER_60_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16346_ _16346_/CLK _16346_/D vssd1 vssd1 vccd1 vccd1 _16346_/Q sky130_fd_sc_hd__dfxtp_1
X_13558_ _16272_/Q _13565_/C _13443_/X vssd1 vssd1 vccd1 vccd1 _13561_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12509_ _13638_/A vssd1 vssd1 vccd1 vccd1 _12739_/B sky130_fd_sc_hd__clkbuf_2
X_16277_ _16346_/CLK _16277_/D vssd1 vssd1 vccd1 vccd1 _16277_/Q sky130_fd_sc_hd__dfxtp_1
X_13489_ _13526_/A _13489_/B _13489_/C vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__and3_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15228_ _15241_/C vssd1 vssd1 vccd1 vccd1 _15248_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15159_ _15180_/A _15159_/B _15163_/B vssd1 vssd1 vccd1 vccd1 _16511_/D sky130_fd_sc_hd__nor3_1
XFILLER_126_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07981_ _16575_/Q _16573_/Q vssd1 vssd1 vccd1 vccd1 _07982_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09720_ _15683_/Q _09867_/B _09727_/C vssd1 vssd1 vccd1 vccd1 _09722_/C sky130_fd_sc_hd__nand3_1
XFILLER_101_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09651_ _09750_/A vssd1 vssd1 vccd1 vccd1 _09651_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08602_ _09815_/A vssd1 vssd1 vccd1 vccd1 _10294_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09582_ _09595_/A _09582_/B _09587_/A vssd1 vssd1 vccd1 vccd1 _15652_/D sky130_fd_sc_hd__nor3_1
XFILLER_82_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08533_ _08521_/A _08521_/B _08532_/X vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__a21o_1
X_08464_ _08399_/A _08399_/B _08463_/Y vssd1 vssd1 vccd1 vccd1 _08466_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08395_ _08395_/A _08395_/B vssd1 vssd1 vccd1 vccd1 _08463_/A sky130_fd_sc_hd__xnor2_4
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09016_ _15540_/Q _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09018_/C sky130_fd_sc_hd__nand3_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09918_ _15721_/Q _09925_/C _09683_/X vssd1 vssd1 vccd1 vccd1 _09921_/A sky130_fd_sc_hd__a21oi_1
XFILLER_59_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09849_ _09849_/A _09849_/B vssd1 vssd1 vccd1 vccd1 _09849_/X sky130_fd_sc_hd__or2_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12860_ _16173_/Q _13082_/B _12860_/C vssd1 vssd1 vccd1 vccd1 _12868_/B sky130_fd_sc_hd__and3_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11811_ _11832_/A _11811_/B _11811_/C vssd1 vssd1 vccd1 vccd1 _11812_/A sky130_fd_sc_hd__and3_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _13638_/A vssd1 vssd1 vccd1 vccd1 _13022_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14814_/A vssd1 vssd1 vccd1 vccd1 _14756_/B sky130_fd_sc_hd__buf_2
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11764_/C vssd1 vssd1 vccd1 vccd1 _11779_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14461_ _14476_/A _14461_/B _14461_/C vssd1 vssd1 vccd1 vccd1 _14462_/A sky130_fd_sc_hd__and3_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11679_/C sky130_fd_sc_hd__nor2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _16555_/Q _16200_/D vssd1 vssd1 vccd1 vccd1 _16200_/Q sky130_fd_sc_hd__dfxtp_1
X_13412_ _13412_/A _13412_/B _13412_/C vssd1 vssd1 vccd1 vccd1 _13413_/A sky130_fd_sc_hd__and3_1
X_10624_ _15839_/Q _15838_/Q _15837_/Q _10476_/X vssd1 vssd1 vccd1 vccd1 _15849_/D
+ sky130_fd_sc_hd__o31a_1
X_14392_ _16460_/Q vssd1 vssd1 vccd1 vccd1 _14406_/C sky130_fd_sc_hd__inv_2
XFILLER_139_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16131_ _16554_/Q _16131_/D vssd1 vssd1 vccd1 vccd1 _16131_/Q sky130_fd_sc_hd__dfxtp_1
X_13343_ _14186_/A vssd1 vssd1 vccd1 vccd1 _13573_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10555_ _10553_/Y _10549_/C _10551_/Y _10552_/X vssd1 vssd1 vccd1 vccd1 _10556_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_139_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16062_ _16118_/CLK _16062_/D vssd1 vssd1 vccd1 vccd1 _16062_/Q sky130_fd_sc_hd__dfxtp_2
X_13274_ _16231_/Q _13383_/B _13283_/C vssd1 vssd1 vccd1 vccd1 _13279_/A sky130_fd_sc_hd__and3_1
X_10486_ _10486_/A vssd1 vssd1 vccd1 vccd1 _10679_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15013_ _15013_/A vssd1 vssd1 vccd1 vccd1 _15027_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12225_ _12225_/A vssd1 vssd1 vccd1 vccd1 _12456_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_12156_ _12156_/A vssd1 vssd1 vccd1 vccd1 _16072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11107_ _11334_/A vssd1 vssd1 vccd1 vccd1 _11148_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12087_ _16064_/Q _12318_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12089_/C sky130_fd_sc_hd__nand3_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11038_ _15916_/Q _11045_/C _10866_/X vssd1 vssd1 vccd1 vccd1 _11038_/Y sky130_fd_sc_hd__a21oi_1
X_15915_ _15365_/A _15915_/D vssd1 vssd1 vccd1 vccd1 _15915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15846_ _16570_/CLK _15846_/D vssd1 vssd1 vccd1 vccd1 _15846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15777_ _15812_/CLK _15777_/D vssd1 vssd1 vccd1 vccd1 _15777_/Q sky130_fd_sc_hd__dfxtp_1
X_12989_ _13009_/C vssd1 vssd1 vccd1 vccd1 _13022_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14728_ _16534_/Q vssd1 vssd1 vccd1 vccd1 _14742_/C sky130_fd_sc_hd__inv_2
XFILLER_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14659_ _14657_/Y _14651_/C _14654_/Y _14664_/A vssd1 vssd1 vccd1 vccd1 _14664_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08180_ _08004_/A _08004_/B _08003_/A vssd1 vssd1 vccd1 vccd1 _08360_/B sky130_fd_sc_hd__o21ai_2
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16329_ _16346_/CLK _16329_/D vssd1 vssd1 vccd1 vccd1 _16329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07964_ _12307_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07965_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09703_ _09658_/X _09701_/B _09651_/X vssd1 vssd1 vccd1 vccd1 _09703_/Y sky130_fd_sc_hd__a21oi_1
X_07895_ _09905_/C _08140_/B vssd1 vssd1 vccd1 vccd1 _07896_/B sky130_fd_sc_hd__xnor2_1
XFILLER_68_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09634_ _09634_/A vssd1 vssd1 vccd1 vccd1 _15662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09565_ _09560_/Y _09563_/X _09564_/Y vssd1 vssd1 vccd1 vccd1 _15647_/D sky130_fd_sc_hd__o21a_1
XFILLER_71_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08516_ _08534_/B _08516_/B vssd1 vssd1 vccd1 vccd1 _08532_/B sky130_fd_sc_hd__xnor2_2
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09496_ _15637_/Q _09669_/B _09496_/C vssd1 vssd1 vccd1 vccd1 _09501_/A sky130_fd_sc_hd__and3_1
XFILLER_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08447_ _08365_/A _08365_/B _08364_/A vssd1 vssd1 vccd1 vccd1 _08453_/A sky130_fd_sc_hd__a21o_1
XFILLER_24_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08378_ _08449_/A _08378_/B vssd1 vssd1 vccd1 vccd1 _08379_/B sky130_fd_sc_hd__or2_2
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ _10340_/A vssd1 vssd1 vccd1 vccd1 _10399_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10271_ _10271_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10271_/X sky130_fd_sc_hd__or2_1
XFILLER_105_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _16053_/Q _12232_/B _12010_/C vssd1 vssd1 vccd1 vccd1 _12018_/B sky130_fd_sc_hd__and3_1
XFILLER_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13961_ _13977_/A _13961_/B _13961_/C vssd1 vssd1 vccd1 vccd1 _13962_/A sky130_fd_sc_hd__and3_1
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15700_ _15791_/CLK _15700_/D vssd1 vssd1 vccd1 vccd1 _15700_/Q sky130_fd_sc_hd__dfxtp_1
X_12912_ _12909_/Y _12918_/A _12911_/Y _12907_/C vssd1 vssd1 vccd1 vccd1 _12914_/B
+ sky130_fd_sc_hd__o211a_1
X_13892_ _13927_/A _13892_/B _13896_/A vssd1 vssd1 vccd1 vccd1 _16318_/D sky130_fd_sc_hd__nor3_1
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15631_ _15812_/CLK _15631_/D vssd1 vssd1 vccd1 vccd1 _15631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ _16171_/Q _13068_/B _12852_/C vssd1 vssd1 vccd1 vccd1 _12843_/X sky130_fd_sc_hd__and3_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ _15812_/CLK _15562_/D vssd1 vssd1 vccd1 vccd1 _15562_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12774_/A vssd1 vssd1 vccd1 vccd1 _16160_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14513_/A vssd1 vssd1 vccd1 vccd1 _16408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11725_ _11805_/A _11725_/B _11731_/B vssd1 vssd1 vccd1 vccd1 _16011_/D sky130_fd_sc_hd__nor3_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _16570_/CLK _15493_/D vssd1 vssd1 vccd1 vccd1 _15493_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14444_ _14444_/A vssd1 vssd1 vccd1 vccd1 _14458_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11656_ _11653_/Y _11654_/X _11655_/Y _11651_/C vssd1 vssd1 vccd1 vccd1 _11658_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_80_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10607_ _15846_/Q _10702_/B _10612_/C vssd1 vssd1 vccd1 vccd1 _10607_/Y sky130_fd_sc_hd__nand3_1
X_14375_ _16387_/Q _14598_/B _14380_/C vssd1 vssd1 vccd1 vccd1 _14375_/Y sky130_fd_sc_hd__nand3_1
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11587_ _11585_/Y _11586_/X _11582_/C _11583_/C vssd1 vssd1 vccd1 vccd1 _11589_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_127_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16114_ _16554_/Q _16114_/D vssd1 vssd1 vccd1 vccd1 _16114_/Q sky130_fd_sc_hd__dfxtp_1
X_13326_ _16239_/Q _13364_/C _13216_/X vssd1 vssd1 vccd1 vccd1 _13328_/B sky130_fd_sc_hd__a21oi_1
X_10538_ _15835_/Q _10546_/C _10432_/X vssd1 vssd1 vccd1 vccd1 _10541_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16045_ _16554_/Q _16045_/D vssd1 vssd1 vccd1 vccd1 _16045_/Q sky130_fd_sc_hd__dfxtp_1
X_13257_ _16229_/Q _13364_/B _13257_/C vssd1 vssd1 vccd1 vccd1 _13266_/B sky130_fd_sc_hd__and3_1
XFILLER_143_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10469_ _10469_/A vssd1 vssd1 vccd1 vccd1 _10469_/X sky130_fd_sc_hd__clkbuf_2
X_12208_ _12208_/A vssd1 vssd1 vccd1 vccd1 _16080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13188_ _13185_/Y _13186_/X _13187_/Y _13181_/C vssd1 vssd1 vccd1 vccd1 _13190_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_2_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12139_ _12152_/C vssd1 vssd1 vccd1 vccd1 _12160_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15829_ _16551_/CLK _15829_/D vssd1 vssd1 vccd1 vccd1 _15829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09350_ _09299_/X _09347_/B _09349_/Y vssd1 vssd1 vccd1 vccd1 _15604_/D sky130_fd_sc_hd__o21a_1
X_08301_ _08301_/A _08316_/A vssd1 vssd1 vccd1 vccd1 _08314_/A sky130_fd_sc_hd__xnor2_2
XFILLER_61_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09281_ _09277_/A _09277_/B _09276_/Y _09280_/Y vssd1 vssd1 vccd1 vccd1 _15592_/D
+ sky130_fd_sc_hd__o31a_1
X_08232_ _16588_/Q _08069_/B _08231_/X vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__a21o_2
XFILLER_21_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08163_ _16593_/Q _16591_/Q _07941_/A vssd1 vssd1 vccd1 vccd1 _08165_/B sky130_fd_sc_hd__a21oi_1
XFILLER_146_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08094_ _08094_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08284_/B sky130_fd_sc_hd__xor2_4
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08996_ _08994_/A _08994_/B _08995_/X vssd1 vssd1 vccd1 vccd1 _15529_/D sky130_fd_sc_hd__a21oi_1
X_07947_ _10583_/C _07947_/B vssd1 vssd1 vccd1 vccd1 _07948_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07878_ _16424_/Q _16406_/Q vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__or2_1
X_09617_ _09898_/A vssd1 vssd1 vccd1 vccd1 _09617_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09548_ _09548_/A vssd1 vssd1 vccd1 vccd1 _15644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09479_ _09699_/A vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _11547_/A _11510_/B _11510_/C vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__and3_1
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12490_ _12505_/A _12490_/B _12490_/C vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__and3_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _12292_/A vssd1 vssd1 vccd1 vccd1 _11441_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14160_ _14160_/A vssd1 vssd1 vccd1 vccd1 _14197_/A sky130_fd_sc_hd__clkbuf_2
X_11372_ _11372_/A vssd1 vssd1 vccd1 vccd1 _15962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13111_ _13392_/A vssd1 vssd1 vccd1 vccd1 _13336_/B sky130_fd_sc_hd__clkbuf_2
X_10323_ _10220_/X _10314_/B _10319_/B _10322_/Y vssd1 vssd1 vccd1 vccd1 _15793_/D
+ sky130_fd_sc_hd__o31a_1
X_14091_ _14091_/A vssd1 vssd1 vccd1 vccd1 _16346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13042_ _13076_/C vssd1 vssd1 vccd1 vccd1 _13082_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10254_ _15783_/Q _10446_/B _10261_/C vssd1 vssd1 vccd1 vccd1 _10254_/X sky130_fd_sc_hd__and3_1
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10185_ _10186_/B _10186_/C _10186_/A vssd1 vssd1 vccd1 vccd1 _10187_/B sky130_fd_sc_hd__a21o_1
XFILLER_132_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14993_ _14993_/A vssd1 vssd1 vccd1 vccd1 _16483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16732_ _16732_/A _07838_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
X_13944_ _13958_/C vssd1 vssd1 vccd1 vccd1 _13966_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13875_ _16317_/Q _13929_/B _13875_/C vssd1 vssd1 vccd1 vccd1 _13883_/B sky130_fd_sc_hd__and3_1
XFILLER_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15614_ _15812_/CLK _15614_/D vssd1 vssd1 vccd1 vccd1 _15614_/Q sky130_fd_sc_hd__dfxtp_1
X_12826_ _16169_/Q _12836_/C _12605_/X vssd1 vssd1 vccd1 vccd1 _12826_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16594_ _16595_/CLK _16594_/D vssd1 vssd1 vccd1 vccd1 _16594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15545_ _15791_/CLK _15545_/D vssd1 vssd1 vccd1 vccd1 _15545_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12770_/C vssd1 vssd1 vccd1 vccd1 _12778_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11706_/Y _11701_/C _11703_/Y _11705_/X vssd1 vssd1 vccd1 vccd1 _11709_/C
+ sky130_fd_sc_hd__a211o_1
X_15476_ _16570_/CLK _15476_/D vssd1 vssd1 vccd1 vccd1 _15476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12688_ _12684_/Y _12694_/A _12687_/Y _12681_/C vssd1 vssd1 vccd1 vccd1 _12690_/B
+ sky130_fd_sc_hd__o211a_1
X_14427_ _16396_/Q _14427_/B _14427_/C vssd1 vssd1 vccd1 vccd1 _14435_/A sky130_fd_sc_hd__and3_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _11637_/Y _11638_/X _11634_/C _11635_/C vssd1 vssd1 vccd1 vccd1 _11641_/B
+ sky130_fd_sc_hd__o211ai_1
X_14358_ _16385_/Q _14414_/B _14358_/C vssd1 vssd1 vccd1 vccd1 _14358_/Y sky130_fd_sc_hd__nand3_1
XFILLER_7_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13309_ _13362_/A _13309_/B _13313_/B vssd1 vssd1 vccd1 vccd1 _16235_/D sky130_fd_sc_hd__nor3_1
X_14289_ _16376_/Q _14289_/B _14296_/C vssd1 vssd1 vccd1 vccd1 _14291_/C sky130_fd_sc_hd__nand3_1
X_16028_ _16554_/Q _16028_/D vssd1 vssd1 vccd1 vccd1 _16028_/Q sky130_fd_sc_hd__dfxtp_1
X_08850_ _08851_/B _08851_/C _08851_/A vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__a21o_1
X_07801_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07801_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08781_ _08781_/A _08781_/B vssd1 vssd1 vccd1 vccd1 _08782_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09402_ _09405_/C vssd1 vssd1 vccd1 vccd1 _09416_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_92_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09333_ _15604_/Q _09340_/C _10750_/B vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__a21oi_1
X_09264_ _09400_/A vssd1 vssd1 vccd1 vccd1 _09374_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08215_ _14222_/A _08016_/B _08214_/Y vssd1 vssd1 vccd1 vccd1 _08373_/B sky130_fd_sc_hd__o21bai_4
X_09195_ _09195_/A _09195_/B vssd1 vssd1 vccd1 vccd1 _09196_/B sky130_fd_sc_hd__nor2_1
X_08146_ _08146_/A vssd1 vssd1 vccd1 vccd1 _08146_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08077_ _15013_/A _08247_/B vssd1 vssd1 vccd1 vccd1 _08248_/B sky130_fd_sc_hd__xnor2_2
XFILLER_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16684__89 vssd1 vssd1 vccd1 vccd1 _16684__89/HI _16760_/A sky130_fd_sc_hd__conb_1
X_08979_ _08980_/B _08980_/C _08980_/A vssd1 vssd1 vccd1 vccd1 _08981_/B sky130_fd_sc_hd__a21o_1
XFILLER_102_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11990_ _11998_/A _11990_/B _11990_/C vssd1 vssd1 vccd1 vccd1 _11991_/A sky130_fd_sc_hd__and3_1
XFILLER_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10941_ _10944_/B _10944_/C _09978_/X vssd1 vssd1 vccd1 vccd1 _10945_/B sky130_fd_sc_hd__o21ai_1
XFILLER_84_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13660_ _16607_/Q vssd1 vssd1 vccd1 vccd1 _13676_/C sky130_fd_sc_hd__inv_2
X_10872_ _10954_/A _10872_/B _10880_/B vssd1 vssd1 vccd1 vccd1 _15891_/D sky130_fd_sc_hd__nor3_1
XFILLER_25_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12611_ _12611_/A vssd1 vssd1 vccd1 vccd1 _16136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13591_ _16277_/Q _13592_/C _13421_/X vssd1 vssd1 vccd1 vccd1 _13593_/A sky130_fd_sc_hd__a21oi_1
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15330_ _15335_/C vssd1 vssd1 vccd1 vccd1 _15346_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12542_ _12542_/A vssd1 vssd1 vccd1 vccd1 _16127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15261_ _16530_/Q _15261_/B _15261_/C vssd1 vssd1 vccd1 vccd1 _15269_/A sky130_fd_sc_hd__and3_1
X_12473_ _12473_/A vssd1 vssd1 vccd1 vccd1 _12487_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14212_ _14437_/A _14217_/C vssd1 vssd1 vccd1 vccd1 _14212_/X sky130_fd_sc_hd__or2_1
X_11424_ _11424_/A vssd1 vssd1 vccd1 vccd1 _15969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15192_ _15192_/A vssd1 vssd1 vccd1 vccd1 _16517_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_8 _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14140_/Y _14141_/X _14142_/Y _14138_/C vssd1 vssd1 vccd1 vccd1 _14145_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_125_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11355_ _11349_/C _11350_/C _11352_/Y _11353_/X vssd1 vssd1 vccd1 vccd1 _11356_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ _15793_/Q _10313_/B _10204_/X vssd1 vssd1 vccd1 vccd1 _10306_/Y sky130_fd_sc_hd__a21oi_1
X_14074_ _14068_/C _14069_/C _14071_/Y _14072_/X vssd1 vssd1 vccd1 vccd1 _14075_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ _11286_/A vssd1 vssd1 vccd1 vccd1 _15949_/D sky130_fd_sc_hd__clkbuf_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ _13023_/Y _13019_/C _13021_/Y _13030_/A vssd1 vssd1 vccd1 vccd1 _13030_/B
+ sky130_fd_sc_hd__a211oi_1
X_10237_ _15781_/Q _10247_/C _10181_/X vssd1 vssd1 vccd1 vccd1 _10240_/B sky130_fd_sc_hd__a21o_1
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10168_ _10418_/A vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10099_ _15757_/Q _10307_/C _10099_/C vssd1 vssd1 vccd1 vccd1 _10108_/A sky130_fd_sc_hd__and3_1
X_14976_ _14970_/C _14971_/C _14973_/Y _14974_/X vssd1 vssd1 vccd1 vccd1 _14977_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16715_ _16715_/A _07818_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
X_13927_ _13927_/A _13927_/B _13931_/B vssd1 vssd1 vccd1 vccd1 _16323_/D sky130_fd_sc_hd__nor3_1
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _13856_/Y _13851_/C _13854_/Y _13855_/X vssd1 vssd1 vccd1 vccd1 _13859_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_50_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12809_ _12847_/A _12809_/B _12809_/C vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__and3_1
X_16577_ _16595_/CLK _16577_/D vssd1 vssd1 vccd1 vccd1 _16577_/Q sky130_fd_sc_hd__dfxtp_1
X_13789_ _13789_/A _13789_/B _13789_/C vssd1 vssd1 vccd1 vccd1 _13790_/C sky130_fd_sc_hd__nand3_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15528_ _15791_/CLK _15528_/D vssd1 vssd1 vccd1 vccd1 _15528_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15459_ _16551_/CLK _15459_/D vssd1 vssd1 vccd1 vccd1 _15459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08000_ _08208_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _08002_/B sky130_fd_sc_hd__xor2_1
XFILLER_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09951_ _09951_/A _09951_/B _09951_/C vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__and3_1
XFILLER_98_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08902_ _15514_/Q _08943_/B _08907_/C vssd1 vssd1 vccd1 vccd1 _08909_/A sky130_fd_sc_hd__and3_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _09880_/A _09880_/B _09879_/Y _09881_/Y vssd1 vssd1 vccd1 vccd1 _15709_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _15338_/A vssd1 vssd1 vccd1 vccd1 _08833_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08764_ _15415_/A vssd1 vssd1 vccd1 vccd1 _08940_/A sky130_fd_sc_hd__buf_2
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08695_ _08693_/A _08693_/B _08694_/X vssd1 vssd1 vccd1 vccd1 _15466_/D sky130_fd_sc_hd__a21oi_1
XFILLER_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09316_ _15615_/Q vssd1 vssd1 vccd1 vccd1 _09320_/C sky130_fd_sc_hd__inv_2
X_09247_ _09207_/X _09246_/A _09129_/X vssd1 vssd1 vccd1 vccd1 _09247_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09178_ _15576_/Q _09220_/B _09178_/C vssd1 vssd1 vccd1 vccd1 _09180_/C sky130_fd_sc_hd__nand3_1
XFILLER_135_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08129_ _08129_/A _08129_/B _08129_/C vssd1 vssd1 vccd1 vccd1 _08130_/B sky130_fd_sc_hd__and3_1
XFILLER_119_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11140_ _11148_/A _11140_/B _11140_/C vssd1 vssd1 vccd1 vccd1 _11141_/A sky130_fd_sc_hd__and3_1
XFILLER_122_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11071_ _11069_/Y _11070_/X _11066_/C _11067_/C vssd1 vssd1 vccd1 vccd1 _11073_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_103_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10022_ _10220_/A _09978_/X _10017_/B _08854_/A vssd1 vssd1 vccd1 vccd1 _10023_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14830_ _14830_/A vssd1 vssd1 vccd1 vccd1 _15055_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11973_ _11974_/B _11974_/C _11974_/A vssd1 vssd1 vccd1 vccd1 _11975_/B sky130_fd_sc_hd__a21o_1
X_14761_ _14761_/A vssd1 vssd1 vccd1 vccd1 _16447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16500_ _16607_/CLK _16500_/D vssd1 vssd1 vccd1 vccd1 _16500_/Q sky130_fd_sc_hd__dfxtp_1
X_10924_ _10922_/Y _10917_/C _10920_/Y _10921_/X vssd1 vssd1 vccd1 vccd1 _10925_/C
+ sky130_fd_sc_hd__a211o_1
X_13712_ _13712_/A _13712_/B vssd1 vssd1 vccd1 vccd1 _13717_/C sky130_fd_sc_hd__nor2_1
XFILLER_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14692_ _14707_/A _14692_/B _14692_/C vssd1 vssd1 vccd1 vccd1 _14693_/A sky130_fd_sc_hd__and3_1
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16431_ _16607_/CLK _16431_/D vssd1 vssd1 vccd1 vccd1 _16431_/Q sky130_fd_sc_hd__dfxtp_1
X_10855_ _10864_/A _10855_/B _10855_/C vssd1 vssd1 vccd1 vccd1 _10856_/A sky130_fd_sc_hd__and3_1
X_13643_ _13643_/A _13643_/B _13647_/B vssd1 vssd1 vccd1 vccd1 _16283_/D sky130_fd_sc_hd__nor3_1
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _16389_/CLK _16362_/D vssd1 vssd1 vccd1 vccd1 _16362_/Q sky130_fd_sc_hd__dfxtp_1
X_13574_ _13571_/Y _13572_/X _13573_/Y _13568_/C vssd1 vssd1 vccd1 vccd1 _13576_/B
+ sky130_fd_sc_hd__o211ai_1
X_10786_ _10786_/A vssd1 vssd1 vccd1 vccd1 _15879_/D sky130_fd_sc_hd__clkbuf_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _15311_/A _15311_/B _15312_/Y vssd1 vssd1 vccd1 vccd1 _16539_/D sky130_fd_sc_hd__o21ba_1
X_12525_ _12526_/B _12526_/C _12416_/X vssd1 vssd1 vccd1 vccd1 _12527_/B sky130_fd_sc_hd__o21ai_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16293_ _16346_/CLK _16293_/D vssd1 vssd1 vccd1 vccd1 _16293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ _15258_/A _15244_/B _15244_/C vssd1 vssd1 vccd1 vccd1 _15245_/A sky130_fd_sc_hd__and3_1
X_12456_ _16116_/Q _12456_/B _12456_/C vssd1 vssd1 vccd1 vccd1 _12464_/A sky130_fd_sc_hd__and3_1
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11407_ _11407_/A _11407_/B _11407_/C vssd1 vssd1 vccd1 vccd1 _11408_/C sky130_fd_sc_hd__nand3_1
X_15175_ _15188_/C vssd1 vssd1 vccd1 vccd1 _15195_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12387_ _16105_/Q _12443_/B _12387_/C vssd1 vssd1 vccd1 vccd1 _12387_/Y sky130_fd_sc_hd__nand3_1
XFILLER_125_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14126_ _16353_/Q _14135_/C _14015_/X vssd1 vssd1 vccd1 vccd1 _14126_/Y sky130_fd_sc_hd__a21oi_1
X_11338_ _11338_/A vssd1 vssd1 vccd1 vccd1 _15957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14057_ _14072_/C vssd1 vssd1 vccd1 vccd1 _14079_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11269_ _11269_/A vssd1 vssd1 vccd1 vccd1 _11495_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13008_ _16194_/Q _13059_/B _13009_/C vssd1 vssd1 vccd1 vccd1 _13008_/X sky130_fd_sc_hd__and3_1
XFILLER_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14959_ _16468_/Q _16467_/Q _16466_/Q _14900_/X vssd1 vssd1 vccd1 vccd1 _16478_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08480_ _08480_/A _08480_/B vssd1 vssd1 vccd1 vccd1 _08481_/B sky130_fd_sc_hd__and2_1
XFILLER_63_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09101_ _09101_/A _09101_/B _09101_/C vssd1 vssd1 vccd1 vccd1 _09102_/C sky130_fd_sc_hd__nand3_1
X_09032_ _09074_/A _09032_/B vssd1 vssd1 vccd1 vccd1 _09032_/X sky130_fd_sc_hd__or2_1
XFILLER_136_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09934_ _09307_/X _09932_/B _09894_/X vssd1 vssd1 vccd1 vccd1 _09934_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09865_ _09946_/A _09865_/B _09869_/A vssd1 vssd1 vccd1 vccd1 _15706_/D sky130_fd_sc_hd__nor3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08816_ _08846_/A _08816_/B _08824_/B vssd1 vssd1 vccd1 vccd1 _15492_/D sky130_fd_sc_hd__nor3_1
X_09796_ _15686_/Q _15685_/Q _15684_/Q _09756_/X vssd1 vssd1 vccd1 vccd1 _15696_/D
+ sky130_fd_sc_hd__o31a_1
X_16654__59 vssd1 vssd1 vccd1 vccd1 _16654__59/HI _16730_/A sky130_fd_sc_hd__conb_1
XFILLER_100_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08747_ _08747_/A vssd1 vssd1 vccd1 vccd1 _08748_/A sky130_fd_sc_hd__buf_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _15468_/Q _08807_/B _08678_/C vssd1 vssd1 vccd1 vccd1 _08680_/C sky130_fd_sc_hd__nand3_1
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10638_/Y _10639_/X _10635_/C _10636_/C vssd1 vssd1 vccd1 vccd1 _10642_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_139_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ _10569_/A _10569_/B _10570_/X vssd1 vssd1 vccd1 vccd1 _15837_/D sky130_fd_sc_hd__a21oi_1
X_12310_ _12346_/C vssd1 vssd1 vccd1 vccd1 _12352_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_139_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13290_ _16234_/Q _13292_/C _13289_/X vssd1 vssd1 vccd1 vccd1 _13290_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12241_ _12468_/A vssd1 vssd1 vccd1 vccd1 _12283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12172_ _16076_/Q _12179_/C _12000_/X vssd1 vssd1 vccd1 vccd1 _12172_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ _11123_/A _11123_/B _11123_/C vssd1 vssd1 vccd1 vccd1 _11124_/C sky130_fd_sc_hd__nand3_1
XFILLER_123_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ _15365_/A _15931_/D vssd1 vssd1 vccd1 vccd1 _15931_/Q sky130_fd_sc_hd__dfxtp_1
X_11054_ _11088_/A _11054_/B _11054_/C vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__and3_1
XFILLER_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10005_ _10005_/A _10005_/B vssd1 vssd1 vccd1 vccd1 _10005_/X sky130_fd_sc_hd__or2_1
XFILLER_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15862_ _16570_/CLK _15862_/D vssd1 vssd1 vccd1 vccd1 _15862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14813_ _16457_/Q _14823_/C _14588_/X vssd1 vssd1 vccd1 vccd1 _14813_/Y sky130_fd_sc_hd__a21oi_1
X_15793_ _15812_/CLK _15793_/D vssd1 vssd1 vccd1 vccd1 _15793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14744_ _14738_/C _14739_/C _14741_/Y _14742_/X vssd1 vssd1 vccd1 vccd1 _14745_/C
+ sky130_fd_sc_hd__a211o_1
X_11956_ _11954_/A _11954_/B _11955_/X vssd1 vssd1 vccd1 vccd1 _16044_/D sky130_fd_sc_hd__a21oi_1
XFILLER_17_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10907_ _15897_/Q _11070_/B _10907_/C vssd1 vssd1 vccd1 vccd1 _10907_/X sky130_fd_sc_hd__and3_1
X_14675_ _14675_/A vssd1 vssd1 vccd1 vccd1 _14689_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11887_ _11885_/Y _11881_/C _11883_/Y _11884_/X vssd1 vssd1 vccd1 vccd1 _11888_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater20 _15812_/CLK vssd1 vssd1 vccd1 vccd1 _16570_/CLK sky130_fd_sc_hd__buf_12
X_16414_ input11/X _16414_/D vssd1 vssd1 vccd1 vccd1 _16414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ _10838_/A _10838_/B _10838_/C vssd1 vssd1 vccd1 vccd1 _10839_/C sky130_fd_sc_hd__nand3_1
X_13626_ _13622_/Y _13623_/X _13625_/Y _13620_/C vssd1 vssd1 vccd1 vccd1 _13628_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16345_ _16346_/CLK _16345_/D vssd1 vssd1 vccd1 vccd1 _16345_/Q sky130_fd_sc_hd__dfxtp_1
X_13557_ _13643_/A _13557_/B _13561_/A vssd1 vssd1 vccd1 vccd1 _16270_/D sky130_fd_sc_hd__nor3_1
XFILLER_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10769_ _10791_/C vssd1 vssd1 vccd1 vccd1 _10805_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12508_ input5/X vssd1 vssd1 vccd1 vccd1 _13638_/A sky130_fd_sc_hd__buf_2
XFILLER_146_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13488_ _13717_/A _13488_/B _13488_/C vssd1 vssd1 vccd1 vccd1 _13489_/C sky130_fd_sc_hd__or3_1
X_16276_ _16533_/Q _16276_/D vssd1 vssd1 vccd1 vccd1 _16276_/Q sky130_fd_sc_hd__dfxtp_1
X_15227_ _16406_/Q vssd1 vssd1 vccd1 vccd1 _15241_/C sky130_fd_sc_hd__inv_2
X_12439_ _12439_/A vssd1 vssd1 vccd1 vccd1 _16112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15158_ _15156_/Y _15152_/C _15154_/Y _15163_/A vssd1 vssd1 vccd1 vccd1 _15163_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_114_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14109_ _14110_/B _14110_/C _14108_/X vssd1 vssd1 vccd1 vccd1 _14111_/B sky130_fd_sc_hd__o21ai_1
X_07980_ _16575_/Q _16573_/Q vssd1 vssd1 vccd1 vccd1 _07982_/A sky130_fd_sc_hd__or2_1
X_15089_ _16501_/Q _15247_/B _15090_/C vssd1 vssd1 vccd1 vccd1 _15089_/X sky130_fd_sc_hd__and3_1
XFILLER_113_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ _09648_/X _09650_/B vssd1 vssd1 vccd1 vccd1 _09650_/X sky130_fd_sc_hd__and2b_1
XFILLER_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08601_ _13060_/A vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09581_ _15655_/Q _09669_/B _09581_/C vssd1 vssd1 vccd1 vccd1 _09587_/A sky130_fd_sc_hd__and3_1
XFILLER_83_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08532_ _08532_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _08532_/X sky130_fd_sc_hd__and2_1
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08463_ _08463_/A _08463_/B vssd1 vssd1 vccd1 vccd1 _08463_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08394_ _08394_/A _08394_/B vssd1 vssd1 vccd1 vccd1 _08395_/B sky130_fd_sc_hd__nor2_2
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09015_ _15540_/Q _09016_/C _09014_/X vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__a21o_1
XFILLER_3_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09917_ _09946_/A _09917_/B _09920_/B vssd1 vssd1 vccd1 vccd1 _15717_/D sky130_fd_sc_hd__nor3_1
XFILLER_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09848_ _09848_/A _09848_/B vssd1 vssd1 vccd1 vccd1 _09849_/B sky130_fd_sc_hd__nor2_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09779_ _09777_/A _09777_/B _09776_/Y _09778_/Y vssd1 vssd1 vccd1 vccd1 _15691_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11810_/A _11810_/B _11810_/C vssd1 vssd1 vccd1 vccd1 _11811_/C sky130_fd_sc_hd__nand3_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _16164_/Q _12798_/C _12567_/X vssd1 vssd1 vccd1 vccd1 _12790_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11757_/C vssd1 vssd1 vccd1 vccd1 _11764_/C sky130_fd_sc_hd__clkbuf_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11672_ _12801_/A vssd1 vssd1 vccd1 vccd1 _11901_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14454_/C _14455_/C _14457_/Y _14458_/X vssd1 vssd1 vccd1 vccd1 _14461_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10623_ _10526_/X _10620_/B _10622_/Y vssd1 vssd1 vccd1 vccd1 _15848_/D sky130_fd_sc_hd__o21a_1
X_13411_ _13409_/Y _13404_/C _13406_/Y _13408_/X vssd1 vssd1 vccd1 vccd1 _13412_/C
+ sky130_fd_sc_hd__a211o_1
X_14391_ _14391_/A vssd1 vssd1 vccd1 vccd1 _16389_/D sky130_fd_sc_hd__clkbuf_1
X_16130_ _16554_/Q _16130_/D vssd1 vssd1 vccd1 vccd1 _16130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13342_ _16242_/Q _13342_/B _13344_/C vssd1 vssd1 vccd1 vccd1 _13342_/X sky130_fd_sc_hd__and3_1
X_10554_ _10551_/Y _10552_/X _10553_/Y _10549_/C vssd1 vssd1 vccd1 vccd1 _10556_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_6_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ _16231_/Q _13311_/C _13216_/X vssd1 vssd1 vccd1 vccd1 _13275_/B sky130_fd_sc_hd__a21oi_1
X_16061_ _16554_/Q _16061_/D vssd1 vssd1 vccd1 vccd1 _16061_/Q sky130_fd_sc_hd__dfxtp_1
X_10485_ _15826_/Q _10494_/C _10432_/X vssd1 vssd1 vccd1 vccd1 _10489_/B sky130_fd_sc_hd__a21o_1
X_15012_ _16477_/Q _16476_/Q _16475_/Q _14900_/X vssd1 vssd1 vccd1 vccd1 _16487_/D
+ sky130_fd_sc_hd__o31a_1
X_12224_ _16084_/Q _12232_/C _12000_/X vssd1 vssd1 vccd1 vccd1 _12224_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_142_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12155_ _12170_/A _12155_/B _12155_/C vssd1 vssd1 vccd1 vccd1 _12156_/A sky130_fd_sc_hd__and3_1
XFILLER_123_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11106_ _11957_/A vssd1 vssd1 vccd1 vccd1 _11334_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12086_ _12373_/A vssd1 vssd1 vccd1 vccd1 _12318_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11037_ _11037_/A vssd1 vssd1 vccd1 vccd1 _15914_/D sky130_fd_sc_hd__clkbuf_1
X_15914_ _15365_/A _15914_/D vssd1 vssd1 vccd1 vccd1 _15914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15845_ _16570_/CLK _15845_/D vssd1 vssd1 vccd1 vccd1 _15845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15776_ _15812_/CLK _15776_/D vssd1 vssd1 vccd1 vccd1 _15776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12988_ _13001_/C vssd1 vssd1 vccd1 vccd1 _13009_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14727_ _16432_/Q _16431_/Q _16430_/Q _14615_/X vssd1 vssd1 vccd1 vccd1 _16442_/D
+ sky130_fd_sc_hd__o31a_1
X_11939_ _11937_/Y _11933_/C _11935_/Y _11936_/X vssd1 vssd1 vccd1 vccd1 _11940_/C
+ sky130_fd_sc_hd__a211o_1
X_14658_ _14654_/Y _14664_/A _14657_/Y _14651_/C vssd1 vssd1 vccd1 vccd1 _14660_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13609_ _13643_/A _13609_/B _13613_/A vssd1 vssd1 vccd1 vccd1 _16278_/D sky130_fd_sc_hd__nor3_1
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14589_ _16421_/Q _14597_/C _14588_/X vssd1 vssd1 vccd1 vccd1 _14589_/Y sky130_fd_sc_hd__a21oi_1
X_16328_ _16346_/CLK _16328_/D vssd1 vssd1 vccd1 vccd1 _16328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16259_ _16261_/CLK _16259_/D vssd1 vssd1 vccd1 vccd1 _16259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07963_ _07963_/A _07963_/B vssd1 vssd1 vccd1 vccd1 _07964_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09702_ _09524_/X _09700_/B _09701_/Y vssd1 vssd1 vccd1 vccd1 _15675_/D sky130_fd_sc_hd__o21a_1
XFILLER_68_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07894_ _10379_/C _07894_/B vssd1 vssd1 vccd1 vccd1 _08140_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16624__29 vssd1 vssd1 vccd1 vccd1 _16624__29/HI _16690_/A sky130_fd_sc_hd__conb_1
X_09633_ _09810_/A _09633_/B _09633_/C vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__and3_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09564_ _09560_/Y _09563_/X _09530_/X vssd1 vssd1 vccd1 vccd1 _09564_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ _08515_/A _08515_/B vssd1 vssd1 vccd1 vccd1 _08516_/B sky130_fd_sc_hd__xnor2_4
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09495_ _09801_/A vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ _08446_/A _08494_/A vssd1 vssd1 vccd1 vccd1 _08472_/A sky130_fd_sc_hd__xnor2_4
XFILLER_51_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08377_ _08377_/A _08377_/B _08377_/C vssd1 vssd1 vccd1 vccd1 _08378_/B sky130_fd_sc_hd__and3_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10270_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13960_ _13953_/C _13954_/C _13956_/Y _13958_/X vssd1 vssd1 vccd1 vccd1 _13961_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12911_ _16179_/Q _12911_/B _12916_/C vssd1 vssd1 vccd1 vccd1 _12911_/Y sky130_fd_sc_hd__nand3_1
XFILLER_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13891_ _16319_/Q _13948_/B _13900_/C vssd1 vssd1 vccd1 vccd1 _13896_/A sky130_fd_sc_hd__and3_1
XFILLER_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15630_ _15812_/CLK _15630_/D vssd1 vssd1 vccd1 vccd1 _15630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _13407_/A vssd1 vssd1 vccd1 vccd1 _13068_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _16551_/CLK _15561_/D vssd1 vssd1 vccd1 vccd1 _15561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12788_/A _12773_/B _12773_/C vssd1 vssd1 vccd1 vccd1 _12774_/A sky130_fd_sc_hd__and3_1
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14535_/A _14512_/B _14512_/C vssd1 vssd1 vccd1 vccd1 _14513_/A sky130_fd_sc_hd__and3_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11722_/Y _11717_/C _11720_/Y _11731_/A vssd1 vssd1 vccd1 vccd1 _11731_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _16570_/CLK _15492_/D vssd1 vssd1 vccd1 vccd1 _15492_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _16002_/Q _11773_/B _11662_/C vssd1 vssd1 vccd1 vccd1 _11655_/Y sky130_fd_sc_hd__nand3_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14443_ _14443_/A vssd1 vssd1 vccd1 vccd1 _16397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _15847_/Q _10652_/B _10606_/C vssd1 vssd1 vccd1 vccd1 _10614_/A sky130_fd_sc_hd__and3_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11586_ _15993_/Q _11638_/B _11586_/C vssd1 vssd1 vccd1 vccd1 _11586_/X sky130_fd_sc_hd__and3_1
X_14374_ _14941_/A vssd1 vssd1 vccd1 vccd1 _14598_/B sky130_fd_sc_hd__clkbuf_2
X_16113_ _16554_/Q _16113_/D vssd1 vssd1 vccd1 vccd1 _16113_/Q sky130_fd_sc_hd__dfxtp_1
X_10537_ _10563_/A _10537_/B _10541_/A vssd1 vssd1 vccd1 vccd1 _15832_/D sky130_fd_sc_hd__nor3_1
XFILLER_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13325_ _13358_/C vssd1 vssd1 vccd1 vccd1 _13364_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16044_ _16554_/Q _16044_/D vssd1 vssd1 vccd1 vccd1 _16044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10468_ _10466_/A _10466_/B _10467_/X vssd1 vssd1 vccd1 vccd1 _15819_/D sky130_fd_sc_hd__a21oi_1
X_13256_ _16229_/Q _13257_/C _13140_/X vssd1 vssd1 vccd1 vccd1 _13258_/A sky130_fd_sc_hd__a21oi_1
X_12207_ _12222_/A _12207_/B _12207_/C vssd1 vssd1 vccd1 vccd1 _12208_/A sky130_fd_sc_hd__and3_1
X_13187_ _16218_/Q _13187_/B _13193_/C vssd1 vssd1 vccd1 vccd1 _13187_/Y sky130_fd_sc_hd__nand3_1
X_10399_ _10399_/A _10399_/B _10399_/C vssd1 vssd1 vccd1 vccd1 _10400_/A sky130_fd_sc_hd__and3_1
XFILLER_124_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12138_ _16580_/Q vssd1 vssd1 vccd1 vccd1 _12152_/C sky130_fd_sc_hd__inv_2
XFILLER_96_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12069_ _12183_/A _12074_/C vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__or2_1
XFILLER_111_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15828_ _16551_/CLK _15828_/D vssd1 vssd1 vccd1 vccd1 _15828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15759_ _15812_/CLK _15759_/D vssd1 vssd1 vccd1 vccd1 _15759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08300_ _08300_/A _08300_/B vssd1 vssd1 vccd1 vccd1 _08316_/A sky130_fd_sc_hd__nand2_1
X_09280_ _09277_/X _09276_/Y _10017_/A vssd1 vssd1 vccd1 vccd1 _09280_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08231_ _16590_/Q _08231_/B vssd1 vssd1 vccd1 vccd1 _08231_/X sky130_fd_sc_hd__and2_1
X_08162_ _12646_/A _07958_/B _07957_/B vssd1 vssd1 vccd1 vccd1 _08165_/A sky130_fd_sc_hd__o21a_2
XFILLER_118_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08093_ _15804_/Q _08280_/B vssd1 vssd1 vccd1 vccd1 _08094_/B sky130_fd_sc_hd__xnor2_2
XFILLER_146_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08995_ _09074_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08995_/X sky130_fd_sc_hd__or2_1
XFILLER_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07946_ _10583_/C _07947_/B vssd1 vssd1 vccd1 vccd1 _07948_/A sky130_fd_sc_hd__or2_1
XFILLER_29_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ _07877_/A _07877_/B vssd1 vssd1 vccd1 vccd1 _07892_/A sky130_fd_sc_hd__or2_4
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09616_ _09615_/X _09611_/B _09572_/X vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__a21oi_1
XFILLER_44_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09547_ _09588_/A _09547_/B _09547_/C vssd1 vssd1 vccd1 vccd1 _09548_/A sky130_fd_sc_hd__and3_1
XFILLER_24_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _09698_/A vssd1 vssd1 vccd1 vccd1 _09656_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08429_ _08414_/A _08414_/B _08428_/X vssd1 vssd1 vccd1 vccd1 _08481_/A sky130_fd_sc_hd__a21oi_1
XFILLER_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11440_ _11520_/A _11440_/B _11446_/B vssd1 vssd1 vccd1 vccd1 _15971_/D sky130_fd_sc_hd__nor3_1
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11371_ _11371_/A _11371_/B _11371_/C vssd1 vssd1 vccd1 vccd1 _11372_/A sky130_fd_sc_hd__and3_1
XFILLER_109_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10322_ _10322_/A _10322_/B vssd1 vssd1 vccd1 vccd1 _10322_/Y sky130_fd_sc_hd__nor2_1
X_13110_ _16209_/Q _13120_/C _12887_/X vssd1 vssd1 vccd1 vccd1 _13110_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14090_ _14090_/A _14090_/B _14090_/C vssd1 vssd1 vccd1 vccd1 _14091_/A sky130_fd_sc_hd__and3_1
XFILLER_124_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041_ _13062_/C vssd1 vssd1 vccd1 vccd1 _13076_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10253_ _15783_/Q _10261_/C _10138_/X vssd1 vssd1 vccd1 vccd1 _10253_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10184_ _15772_/Q _10434_/B _10190_/C vssd1 vssd1 vccd1 vccd1 _10186_/C sky130_fd_sc_hd__nand3_1
XFILLER_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14992_ _14992_/A _14992_/B _14992_/C vssd1 vssd1 vccd1 vccd1 _14993_/A sky130_fd_sc_hd__and3_1
XFILLER_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16731_ _16731_/A _07836_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13943_ _13943_/A vssd1 vssd1 vccd1 vccd1 _13958_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13874_ _16317_/Q _13875_/C _13705_/X vssd1 vssd1 vccd1 vccd1 _13876_/A sky130_fd_sc_hd__a21oi_1
XFILLER_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15613_ _15812_/CLK _15613_/D vssd1 vssd1 vccd1 vccd1 _15613_/Q sky130_fd_sc_hd__dfxtp_1
X_12825_ _12825_/A vssd1 vssd1 vccd1 vccd1 _16167_/D sky130_fd_sc_hd__clkbuf_1
X_16593_ _16595_/CLK _16593_/D vssd1 vssd1 vccd1 vccd1 _16593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15544_ _15791_/CLK _15544_/D vssd1 vssd1 vccd1 vccd1 _15544_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _16591_/Q vssd1 vssd1 vccd1 vccd1 _12770_/C sky130_fd_sc_hd__inv_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11703_/Y _11705_/X _11706_/Y _11701_/C vssd1 vssd1 vccd1 vccd1 _11709_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _16551_/CLK _15475_/D vssd1 vssd1 vccd1 vccd1 _15475_/Q sky130_fd_sc_hd__dfxtp_2
X_12687_ _16147_/Q _12911_/B _12692_/C vssd1 vssd1 vccd1 vccd1 _12687_/Y sky130_fd_sc_hd__nand3_1
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14426_ _16396_/Q _14433_/C _14258_/X vssd1 vssd1 vccd1 vccd1 _14426_/Y sky130_fd_sc_hd__a21oi_1
X_11638_ _16001_/Q _11638_/B _11638_/C vssd1 vssd1 vccd1 vccd1 _11638_/X sky130_fd_sc_hd__and3_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14357_ _16386_/Q _14464_/B _14358_/C vssd1 vssd1 vccd1 vccd1 _14357_/X sky130_fd_sc_hd__and3_1
XFILLER_116_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11569_ _11737_/A _11569_/B _11569_/C vssd1 vssd1 vccd1 vccd1 _11570_/C sky130_fd_sc_hd__or3_1
X_13308_ _13306_/Y _13302_/C _13304_/Y _13313_/A vssd1 vssd1 vccd1 vccd1 _13313_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14288_ _16376_/Q _14296_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14291_/B sky130_fd_sc_hd__a21o_1
X_16027_ _16554_/Q _16027_/D vssd1 vssd1 vccd1 vccd1 _16027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13239_ _13239_/A vssd1 vssd1 vccd1 vccd1 _16225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07800_ _07806_/A vssd1 vssd1 vccd1 vccd1 _07805_/A sky130_fd_sc_hd__buf_6
X_08780_ _08780_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08782_/A sky130_fd_sc_hd__or2_1
XFILLER_111_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09401_ _15633_/Q vssd1 vssd1 vccd1 vccd1 _09405_/C sky130_fd_sc_hd__inv_2
XFILLER_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09332_ _09374_/A _09332_/B _09335_/B vssd1 vssd1 vccd1 vccd1 _15600_/D sky130_fd_sc_hd__nor3_1
XFILLER_34_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09263_ _09263_/A vssd1 vssd1 vccd1 vccd1 _15590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08214_ _14335_/A _08214_/B vssd1 vssd1 vccd1 vccd1 _08214_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ _09194_/A _09194_/B vssd1 vssd1 vccd1 vccd1 _09195_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08145_ _08145_/A _08319_/A vssd1 vssd1 vccd1 vccd1 _08291_/A sky130_fd_sc_hd__xnor2_1
XFILLER_107_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08076_ _08256_/A _08076_/B vssd1 vssd1 vccd1 vccd1 _08247_/B sky130_fd_sc_hd__xnor2_4
XFILLER_146_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08978_ _15531_/Q _09016_/B _08978_/C vssd1 vssd1 vccd1 vccd1 _08980_/C sky130_fd_sc_hd__nand3_1
XFILLER_69_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07929_ _13269_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _07930_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10940_ _11051_/A vssd1 vssd1 vccd1 vccd1 _10981_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10871_ _10869_/Y _10864_/C _10867_/Y _10880_/A vssd1 vssd1 vccd1 vccd1 _10880_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _12625_/A _12610_/B _12610_/C vssd1 vssd1 vccd1 vccd1 _12611_/A sky130_fd_sc_hd__and3_1
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13590_ _13643_/A _13590_/B _13594_/B vssd1 vssd1 vccd1 vccd1 _16275_/D sky130_fd_sc_hd__nor3_1
XFILLER_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12541_ _12565_/A _12541_/B _12541_/C vssd1 vssd1 vccd1 vccd1 _12542_/A sky130_fd_sc_hd__and3_1
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15260_ _16530_/Q _15267_/C _08747_/A vssd1 vssd1 vccd1 vccd1 _15260_/Y sky130_fd_sc_hd__a21oi_1
X_12472_ _12472_/A vssd1 vssd1 vccd1 vccd1 _16117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14211_ _14211_/A _14211_/B vssd1 vssd1 vccd1 vccd1 _14217_/C sky130_fd_sc_hd__nor2_1
XFILLER_138_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11423_ _11431_/A _11423_/B _11423_/C vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__and3_1
X_15191_ _15205_/A _15191_/B _15191_/C vssd1 vssd1 vccd1 vccd1 _15192_/A sky130_fd_sc_hd__and3_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_9 _14906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11354_ _11352_/Y _11353_/X _11349_/C _11350_/C vssd1 vssd1 vccd1 vccd1 _11356_/B
+ sky130_fd_sc_hd__o211ai_1
X_14142_ _16354_/Q _14311_/B _14148_/C vssd1 vssd1 vccd1 vccd1 _14142_/Y sky130_fd_sc_hd__nand3_1
XFILLER_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ _10305_/A vssd1 vssd1 vccd1 vccd1 _15790_/D sky130_fd_sc_hd__clkbuf_1
X_11285_ _11319_/A _11285_/B _11285_/C vssd1 vssd1 vccd1 vccd1 _11286_/A sky130_fd_sc_hd__and3_1
X_14073_ _14071_/Y _14072_/X _14068_/C _14069_/C vssd1 vssd1 vccd1 vccd1 _14075_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10236_ _10311_/A _10236_/B _10240_/A vssd1 vssd1 vccd1 vccd1 _15778_/D sky130_fd_sc_hd__nor3_1
X_13024_ _13021_/Y _13030_/A _13023_/Y _13019_/C vssd1 vssd1 vccd1 vccd1 _13026_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10167_ _09851_/X _10159_/B _10162_/B _10166_/Y vssd1 vssd1 vccd1 vccd1 _15766_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10098_ _15757_/Q _10106_/C _10009_/B vssd1 vssd1 vccd1 vccd1 _10098_/Y sky130_fd_sc_hd__a21oi_1
X_14975_ _14973_/Y _14974_/X _14970_/C _14971_/C vssd1 vssd1 vccd1 vccd1 _14977_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16714_ _16714_/A _07817_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13926_ _13924_/Y _13918_/C _13920_/Y _13931_/A vssd1 vssd1 vccd1 vccd1 _13931_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13857_ _13854_/Y _13855_/X _13856_/Y _13851_/C vssd1 vssd1 vccd1 vccd1 _13859_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ _12868_/A _12808_/B _12808_/C vssd1 vssd1 vccd1 vccd1 _12809_/C sky130_fd_sc_hd__or3_1
X_16576_ _16595_/CLK _16576_/D vssd1 vssd1 vccd1 vccd1 _16576_/Q sky130_fd_sc_hd__dfxtp_1
X_13788_ _13789_/B _13789_/C _13789_/A vssd1 vssd1 vccd1 vccd1 _13790_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15527_ _15791_/CLK _15527_/D vssd1 vssd1 vccd1 vccd1 _15527_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _16156_/Q _12739_/B _12739_/C vssd1 vssd1 vccd1 vccd1 _12747_/A sky130_fd_sc_hd__and3_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ _16551_/CLK _15458_/D vssd1 vssd1 vccd1 vccd1 _15458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14409_ _14424_/A _14409_/B _14409_/C vssd1 vssd1 vccd1 vccd1 _14410_/A sky130_fd_sc_hd__and3_1
XFILLER_129_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15389_ _16021_/Q _16020_/Q _16019_/Q _15385_/X vssd1 vssd1 vccd1 vccd1 _16573_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_128_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09950_ _09950_/A _09950_/B _09950_/C vssd1 vssd1 vccd1 vccd1 _09951_/C sky130_fd_sc_hd__nand3_1
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08901_ _15514_/Q _08907_/C _08859_/X vssd1 vssd1 vccd1 vccd1 _08901_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09880_/X _09879_/Y _09644_/X vssd1 vssd1 vccd1 vccd1 _09881_/Y sky130_fd_sc_hd__a21oi_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _09038_/A vssd1 vssd1 vccd1 vccd1 _08832_/X sky130_fd_sc_hd__clkbuf_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _13652_/A vssd1 vssd1 vccd1 vccd1 _15415_/A sky130_fd_sc_hd__buf_8
XFILLER_26_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08694_ _08870_/A _08694_/B vssd1 vssd1 vccd1 vccd1 _08694_/X sky130_fd_sc_hd__or2_1
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09315_ _15587_/Q _15586_/Q _15585_/Q _09314_/X vssd1 vssd1 vccd1 vccd1 _15597_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_22_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _09246_/A _09246_/B vssd1 vssd1 vccd1 vccd1 _15586_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ _15576_/Q _09178_/C _09014_/X vssd1 vssd1 vccd1 vccd1 _09180_/B sky130_fd_sc_hd__a21o_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ _08129_/A _08129_/B _08129_/C vssd1 vssd1 vccd1 vccd1 _08343_/A sky130_fd_sc_hd__a21oi_4
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08059_ _09761_/C _08059_/B vssd1 vssd1 vccd1 vccd1 _08245_/A sky130_fd_sc_hd__xnor2_4
XFILLER_150_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11070_ _15921_/Q _11070_/B _11070_/C vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__and3_1
XFILLER_150_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10021_ _08654_/X _10017_/B _09792_/X vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__a21oi_1
XFILLER_1_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14760_ _14760_/A _14760_/B _14760_/C vssd1 vssd1 vccd1 vccd1 _14761_/A sky130_fd_sc_hd__and3_1
X_11972_ _16048_/Q _12031_/B _11979_/C vssd1 vssd1 vccd1 vccd1 _11974_/C sky130_fd_sc_hd__nand3_1
X_13711_ _13711_/A _13711_/B vssd1 vssd1 vccd1 vccd1 _13712_/B sky130_fd_sc_hd__nor2_1
X_10923_ _10920_/Y _10921_/X _10922_/Y _10917_/C vssd1 vssd1 vccd1 vccd1 _10925_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14691_ _14685_/C _14686_/C _14688_/Y _14689_/X vssd1 vssd1 vccd1 vccd1 _14692_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16430_ _16607_/CLK _16430_/D vssd1 vssd1 vccd1 vccd1 _16430_/Q sky130_fd_sc_hd__dfxtp_1
X_13642_ _13640_/Y _13635_/C _13637_/Y _13647_/A vssd1 vssd1 vccd1 vccd1 _13647_/B
+ sky130_fd_sc_hd__a211oi_1
X_10854_ _10852_/Y _10847_/C _10849_/Y _10851_/X vssd1 vssd1 vccd1 vccd1 _10855_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_25_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16389_/CLK _16361_/D vssd1 vssd1 vccd1 vccd1 _16361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _16273_/Q _13573_/B _13573_/C vssd1 vssd1 vccd1 vccd1 _13573_/Y sky130_fd_sc_hd__nand3_1
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10785_ _10801_/A _10785_/B _10785_/C vssd1 vssd1 vccd1 vccd1 _10786_/A sky130_fd_sc_hd__and3_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15312_/A _15312_/B vssd1 vssd1 vccd1 vccd1 _15312_/Y sky130_fd_sc_hd__nand2_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _12751_/A vssd1 vssd1 vccd1 vccd1 _12565_/A sky130_fd_sc_hd__clkbuf_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _16346_/CLK _16292_/D vssd1 vssd1 vccd1 vccd1 _16292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15243_ _15237_/C _15238_/C _15240_/Y _15241_/X vssd1 vssd1 vccd1 vccd1 _15244_/C
+ sky130_fd_sc_hd__a211o_1
X_12455_ _16116_/Q _12462_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12455_/Y sky130_fd_sc_hd__a21oi_1
X_11406_ _11407_/B _11407_/C _11407_/A vssd1 vssd1 vccd1 vccd1 _11408_/B sky130_fd_sc_hd__a21o_1
XFILLER_138_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15174_ _16532_/Q vssd1 vssd1 vccd1 vccd1 _15188_/C sky130_fd_sc_hd__inv_2
X_12386_ _16106_/Q _12493_/B _12387_/C vssd1 vssd1 vccd1 vccd1 _12386_/X sky130_fd_sc_hd__and3_1
XFILLER_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14125_ _14125_/A vssd1 vssd1 vccd1 vccd1 _16351_/D sky130_fd_sc_hd__clkbuf_1
X_11337_ _11371_/A _11337_/B _11337_/C vssd1 vssd1 vccd1 vccd1 _11338_/A sky130_fd_sc_hd__and3_1
XFILLER_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14056_ _16614_/Q vssd1 vssd1 vccd1 vccd1 _14072_/C sky130_fd_sc_hd__inv_2
X_11268_ _15948_/Q _11322_/B _11268_/C vssd1 vssd1 vccd1 vccd1 _11277_/A sky130_fd_sc_hd__and3_1
XFILLER_97_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _16194_/Q _13009_/C _13006_/X vssd1 vssd1 vccd1 vccd1 _13007_/Y sky130_fd_sc_hd__a21oi_1
X_10219_ _10217_/A _10217_/B _10218_/X vssd1 vssd1 vccd1 vccd1 _15774_/D sky130_fd_sc_hd__a21oi_1
X_11199_ _11197_/Y _11193_/C _11195_/Y _11196_/X vssd1 vssd1 vccd1 vccd1 _11200_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_94_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14958_ _14958_/A vssd1 vssd1 vccd1 vccd1 _16477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ _13905_/Y _13906_/X _13908_/Y _13903_/C vssd1 vssd1 vccd1 vccd1 _13911_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14889_ _14889_/A _14889_/B vssd1 vssd1 vccd1 vccd1 _14890_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16559_ _16595_/CLK _16559_/D vssd1 vssd1 vccd1 vccd1 _16559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09100_ _09101_/B _09101_/C _09101_/A vssd1 vssd1 vccd1 vccd1 _09102_/B sky130_fd_sc_hd__a21o_1
X_09031_ _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _09032_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09933_ _09744_/X _09931_/B _09932_/Y vssd1 vssd1 vccd1 vccd1 _15720_/D sky130_fd_sc_hd__o21a_1
XFILLER_89_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09864_ _15709_/Q _09945_/B _09864_/C vssd1 vssd1 vccd1 vccd1 _09869_/A sky130_fd_sc_hd__and3_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08815_ _08809_/C _08810_/C _08812_/Y _08824_/A vssd1 vssd1 vccd1 vccd1 _08824_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09795_ _09795_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _15695_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08746_ _12849_/A vssd1 vssd1 vccd1 vccd1 _08747_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _15468_/Q _08678_/C _15335_/B vssd1 vssd1 vccd1 vccd1 _08680_/B sky130_fd_sc_hd__a21o_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10570_ _10759_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _10570_/X sky130_fd_sc_hd__or2_1
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09229_ _09256_/A _09229_/B _09233_/B vssd1 vssd1 vccd1 vccd1 _15582_/D sky130_fd_sc_hd__nor3_1
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12240_ _13371_/A vssd1 vssd1 vccd1 vccd1 _12468_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ _12171_/A vssd1 vssd1 vccd1 vccd1 _16074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11122_ _11123_/B _11123_/C _11123_/A vssd1 vssd1 vccd1 vccd1 _11124_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15930_ _16005_/CLK _15930_/D vssd1 vssd1 vccd1 vccd1 _15930_/Q sky130_fd_sc_hd__dfxtp_1
X_11053_ _11169_/A _11053_/B _11053_/C vssd1 vssd1 vccd1 vccd1 _11054_/C sky130_fd_sc_hd__or3_1
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10004_ _10004_/A _10004_/B vssd1 vssd1 vccd1 vccd1 _10004_/Y sky130_fd_sc_hd__nor2_1
X_15861_ _16595_/CLK _15861_/D vssd1 vssd1 vccd1 vccd1 _15861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14812_ _14812_/A vssd1 vssd1 vccd1 vccd1 _16455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15792_ _15812_/CLK _15792_/D vssd1 vssd1 vccd1 vccd1 _15792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14743_ _14741_/Y _14742_/X _14738_/C _14739_/C vssd1 vssd1 vccd1 vccd1 _14745_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11955_ _12183_/A _11960_/C vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__or2_1
X_10906_ _15897_/Q _10914_/C _10905_/X vssd1 vssd1 vccd1 vccd1 _10906_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _16423_/Q _16422_/Q _16421_/Q _14615_/X vssd1 vssd1 vccd1 vccd1 _16433_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_72_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11886_ _11883_/Y _11884_/X _11885_/Y _11881_/C vssd1 vssd1 vccd1 vccd1 _11888_/B
+ sky130_fd_sc_hd__o211ai_1
X_16413_ input11/X _16413_/D vssd1 vssd1 vccd1 vccd1 _16413_/Q sky130_fd_sc_hd__dfxtp_1
X_13625_ _16281_/Q _13856_/B _13625_/C vssd1 vssd1 vccd1 vccd1 _13625_/Y sky130_fd_sc_hd__nand3_1
XFILLER_60_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater21 _15812_/CLK vssd1 vssd1 vccd1 vccd1 _15791_/CLK sky130_fd_sc_hd__buf_12
X_10837_ _10838_/B _10838_/C _10838_/A vssd1 vssd1 vccd1 vccd1 _10839_/B sky130_fd_sc_hd__a21o_1
X_16344_ _16389_/CLK _16344_/D vssd1 vssd1 vccd1 vccd1 _16344_/Q sky130_fd_sc_hd__dfxtp_1
X_13556_ _16271_/Q _13665_/B _13565_/C vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__and3_1
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10768_ _10782_/C vssd1 vssd1 vccd1 vccd1 _10791_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12507_ _16124_/Q _12516_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12507_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16275_ _16533_/Q _16275_/D vssd1 vssd1 vccd1 vccd1 _16275_/Q sky130_fd_sc_hd__dfxtp_1
X_13487_ _14331_/A vssd1 vssd1 vccd1 vccd1 _13717_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10699_ _15865_/Q _10707_/C _09604_/A vssd1 vssd1 vccd1 vccd1 _10699_/Y sky130_fd_sc_hd__a21oi_1
X_15226_ _16513_/Q _16512_/Q _16511_/Q _15172_/X vssd1 vssd1 vccd1 vccd1 _16523_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12438_ _12453_/A _12438_/B _12438_/C vssd1 vssd1 vccd1 vccd1 _12439_/A sky130_fd_sc_hd__and3_1
X_15157_ _15154_/Y _15163_/A _15156_/Y _15152_/C vssd1 vssd1 vccd1 vccd1 _15159_/B
+ sky130_fd_sc_hd__o211a_1
X_12369_ _16103_/Q _12409_/C _12368_/X vssd1 vssd1 vccd1 vccd1 _12371_/B sky130_fd_sc_hd__a21oi_1
XFILLER_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14108_ _14669_/A vssd1 vssd1 vccd1 vccd1 _14108_/X sky130_fd_sc_hd__clkbuf_2
X_15088_ _16501_/Q _15090_/C _14979_/X vssd1 vssd1 vccd1 vccd1 _15088_/Y sky130_fd_sc_hd__a21oi_1
X_14039_ _16339_/Q _14039_/B _14044_/C vssd1 vssd1 vccd1 vccd1 _14039_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08600_ _12886_/A vssd1 vssd1 vccd1 vccd1 _13060_/A sky130_fd_sc_hd__buf_6
XFILLER_94_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09580_ _15655_/Q _09603_/C _09493_/X vssd1 vssd1 vccd1 vccd1 _09582_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08531_ _08529_/A _08529_/B _08530_/Y vssd1 vssd1 vccd1 vccd1 _15450_/D sky130_fd_sc_hd__o21ba_1
X_08462_ _08462_/A _08462_/B vssd1 vssd1 vccd1 vccd1 _08466_/A sky130_fd_sc_hd__xnor2_1
X_08393_ _08393_/A _08393_/B vssd1 vssd1 vccd1 vccd1 _08394_/B sky130_fd_sc_hd__and2_1
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09014_ _09056_/A vssd1 vssd1 vccd1 vccd1 _09014_/X sky130_fd_sc_hd__buf_2
XFILLER_145_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09916_ _09910_/C _09911_/C _09913_/Y _09920_/A vssd1 vssd1 vccd1 vccd1 _09920_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09847_ _09847_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__nor2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09778_ _09777_/X _09776_/Y _09644_/X vssd1 vssd1 vccd1 vccd1 _09778_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _08723_/C _08724_/C _08726_/Y _08734_/A vssd1 vssd1 vccd1 vccd1 _08734_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _16573_/Q vssd1 vssd1 vccd1 vccd1 _11757_/C sky130_fd_sc_hd__inv_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _13085_/A vssd1 vssd1 vccd1 vccd1 _12801_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13410_ _13406_/Y _13408_/X _13409_/Y _13404_/C vssd1 vssd1 vccd1 vccd1 _13412_/B
+ sky130_fd_sc_hd__o211ai_1
X_10622_ _10418_/X _10620_/B _10473_/X vssd1 vssd1 vccd1 vccd1 _10622_/Y sky130_fd_sc_hd__a21oi_1
X_14390_ _14424_/A _14390_/B _14390_/C vssd1 vssd1 vccd1 vccd1 _14391_/A sky130_fd_sc_hd__and3_1
XFILLER_139_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13341_ _16242_/Q _13344_/C _13289_/X vssd1 vssd1 vccd1 vccd1 _13341_/Y sky130_fd_sc_hd__a21oi_1
X_10553_ _15836_/Q _10646_/B _10559_/C vssd1 vssd1 vccd1 vccd1 _10553_/Y sky130_fd_sc_hd__nand3_1
XFILLER_139_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16060_ _16554_/Q _16060_/D vssd1 vssd1 vccd1 vccd1 _16060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13272_ _13305_/C vssd1 vssd1 vccd1 vccd1 _13311_/C sky130_fd_sc_hd__clkbuf_2
X_10484_ _10563_/A _10484_/B _10489_/A vssd1 vssd1 vccd1 vccd1 _15823_/D sky130_fd_sc_hd__nor3_1
XFILLER_6_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15011_ _15011_/A vssd1 vssd1 vccd1 vccd1 _16486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12223_ _12223_/A vssd1 vssd1 vccd1 vccd1 _16082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12154_ _12148_/C _12149_/C _12151_/Y _12152_/X vssd1 vssd1 vccd1 vccd1 _12155_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_123_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11105_ _11103_/A _11103_/B _11104_/X vssd1 vssd1 vccd1 vccd1 _15924_/D sky130_fd_sc_hd__a21oi_1
XFILLER_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12085_ _16064_/Q _12093_/C _12029_/X vssd1 vssd1 vccd1 vccd1 _12089_/B sky130_fd_sc_hd__a21o_1
X_11036_ _11036_/A _11036_/B _11036_/C vssd1 vssd1 vccd1 vccd1 _11037_/A sky130_fd_sc_hd__and3_1
X_15913_ _16553_/Q _15913_/D vssd1 vssd1 vccd1 vccd1 _15913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15844_ _16570_/CLK _15844_/D vssd1 vssd1 vccd1 vccd1 _15844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15775_ _15812_/CLK _15775_/D vssd1 vssd1 vccd1 vccd1 _15775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12987_ _12987_/A vssd1 vssd1 vccd1 vccd1 _13001_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14726_ _14726_/A vssd1 vssd1 vccd1 vccd1 _16441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11938_ _11935_/Y _11936_/X _11937_/Y _11933_/C vssd1 vssd1 vccd1 vccd1 _11940_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_33_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14657_ _16430_/Q _14882_/B _14662_/C vssd1 vssd1 vccd1 vccd1 _14657_/Y sky130_fd_sc_hd__nand3_1
X_11869_ _16033_/Q _11922_/B _11869_/C vssd1 vssd1 vccd1 vccd1 _11869_/X sky130_fd_sc_hd__and3_1
X_13608_ _16279_/Q _13665_/B _13617_/C vssd1 vssd1 vccd1 vccd1 _13613_/A sky130_fd_sc_hd__and3_1
X_14588_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14588_/X sky130_fd_sc_hd__clkbuf_4
X_16327_ _16346_/CLK _16327_/D vssd1 vssd1 vccd1 vccd1 _16327_/Q sky130_fd_sc_hd__dfxtp_1
X_13539_ _13539_/A _13548_/B vssd1 vssd1 vccd1 vccd1 _13541_/A sky130_fd_sc_hd__or2_1
XFILLER_146_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16258_ _16261_/CLK _16258_/D vssd1 vssd1 vccd1 vccd1 _16258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15209_ _16521_/Q _15261_/B _15209_/C vssd1 vssd1 vccd1 vccd1 _15217_/A sky130_fd_sc_hd__and3_1
X_16189_ _16555_/Q _16189_/D vssd1 vssd1 vccd1 vccd1 _16189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07962_ _16581_/Q _16579_/Q vssd1 vssd1 vccd1 vccd1 _07963_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09701_ _09932_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _09701_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07893_ _15840_/Q _08121_/B vssd1 vssd1 vccd1 vccd1 _07894_/B sky130_fd_sc_hd__xnor2_1
X_09632_ _09632_/A _09632_/B _09632_/C vssd1 vssd1 vccd1 vccd1 _09633_/C sky130_fd_sc_hd__nand3_1
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09563_ _09561_/X _09563_/B vssd1 vssd1 vccd1 vccd1 _09563_/X sky130_fd_sc_hd__and2b_1
XFILLER_82_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08514_ _08535_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _08515_/B sky130_fd_sc_hd__xor2_4
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09494_ _15637_/Q _09519_/C _09493_/X vssd1 vssd1 vccd1 vccd1 _09497_/B sky130_fd_sc_hd__a21oi_1
XFILLER_130_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08445_ _08445_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08494_/A sky130_fd_sc_hd__xnor2_2
XFILLER_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ _08377_/A _08377_/B _08377_/C vssd1 vssd1 vccd1 vccd1 _08449_/A sky130_fd_sc_hd__a21oi_1
XFILLER_149_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12910_ _16180_/Q _13022_/B _12910_/C vssd1 vssd1 vccd1 vccd1 _12918_/A sky130_fd_sc_hd__and3_1
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ _16319_/Q _13929_/C _13781_/X vssd1 vssd1 vccd1 vccd1 _13892_/B sky130_fd_sc_hd__a21oi_1
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ _16171_/Q _12852_/C _12619_/X vssd1 vssd1 vccd1 vccd1 _12841_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _16551_/CLK _15560_/D vssd1 vssd1 vccd1 vccd1 _15560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12766_/C _12767_/C _12769_/Y _12770_/X vssd1 vssd1 vccd1 vccd1 _12773_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14511_/A _14511_/B _14511_/C vssd1 vssd1 vccd1 vccd1 _14512_/C sky130_fd_sc_hd__nand3_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11720_/Y _11731_/A _11722_/Y _11717_/C vssd1 vssd1 vccd1 vccd1 _11725_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _16570_/CLK _15491_/D vssd1 vssd1 vccd1 vccd1 _15491_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14476_/A _14442_/B _14442_/C vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__and3_1
X_11654_ _16003_/Q _11654_/B _11662_/C vssd1 vssd1 vccd1 vccd1 _11654_/X sky130_fd_sc_hd__and3_1
XFILLER_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10605_ _15847_/Q _10612_/C _10454_/X vssd1 vssd1 vccd1 vccd1 _10605_/Y sky130_fd_sc_hd__a21oi_1
X_14373_ _16388_/Q _14427_/B _14373_/C vssd1 vssd1 vccd1 vccd1 _14382_/A sky130_fd_sc_hd__and3_1
X_11585_ _15993_/Q _11594_/C _11471_/X vssd1 vssd1 vccd1 vccd1 _11585_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16112_ _16554_/Q _16112_/D vssd1 vssd1 vccd1 vccd1 _16112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13324_ _13344_/C vssd1 vssd1 vccd1 vccd1 _13358_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10536_ _15834_/Q _10726_/B _10536_/C vssd1 vssd1 vccd1 vccd1 _10541_/A sky130_fd_sc_hd__and3_1
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16043_ _16118_/CLK _16043_/D vssd1 vssd1 vccd1 vccd1 _16043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13255_ _13362_/A _13255_/B _13259_/B vssd1 vssd1 vccd1 vccd1 _16227_/D sky130_fd_sc_hd__nor3_1
XFILLER_50_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _10521_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__or2_1
XFILLER_136_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12206_ _12200_/C _12201_/C _12203_/Y _12204_/X vssd1 vssd1 vccd1 vccd1 _12207_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_142_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _16219_/Q _13350_/B _13193_/C vssd1 vssd1 vccd1 vccd1 _13186_/X sky130_fd_sc_hd__and3_1
X_10398_ _10396_/Y _10391_/C _10394_/Y _10395_/X vssd1 vssd1 vccd1 vccd1 _10399_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12137_ _12137_/A vssd1 vssd1 vccd1 vccd1 _16069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12068_ _12068_/A _12068_/B vssd1 vssd1 vccd1 vccd1 _12074_/C sky130_fd_sc_hd__nor2_1
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ _11017_/Y _11018_/X _11014_/C _11015_/C vssd1 vssd1 vccd1 vccd1 _11021_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15827_ _16570_/CLK _15827_/D vssd1 vssd1 vccd1 vccd1 _15827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15758_ _15812_/CLK _15758_/D vssd1 vssd1 vccd1 vccd1 _15758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14709_ _16440_/Q _14716_/C _14537_/X vssd1 vssd1 vccd1 vccd1 _14709_/Y sky130_fd_sc_hd__a21oi_1
X_15689_ _15791_/CLK _15689_/D vssd1 vssd1 vccd1 vccd1 _15689_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08230_ _08051_/A _08228_/Y _08229_/Y vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__a21o_1
XFILLER_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08161_ _13269_/A _07929_/B _07928_/B vssd1 vssd1 vccd1 vccd1 _08171_/A sky130_fd_sc_hd__o21a_1
XFILLER_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08092_ _08092_/A _08092_/B vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__xor2_2
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08994_ _08994_/A _08994_/B vssd1 vssd1 vccd1 vccd1 _08995_/B sky130_fd_sc_hd__nor2_1
XFILLER_102_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07945_ _07945_/A _07945_/B vssd1 vssd1 vccd1 vccd1 _07947_/B sky130_fd_sc_hd__xor2_4
XFILLER_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07876_ _12928_/A _07876_/B vssd1 vssd1 vccd1 vccd1 _07877_/B sky130_fd_sc_hd__and2_1
XFILLER_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09615_ _09615_/A vssd1 vssd1 vccd1 vccd1 _09615_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ _09546_/A _09546_/B _09546_/C vssd1 vssd1 vccd1 vccd1 _09547_/C sky130_fd_sc_hd__nand3_1
XFILLER_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09477_ _09471_/Y _09472_/X _09474_/B vssd1 vssd1 vccd1 vccd1 _09480_/B sky130_fd_sc_hd__o21a_1
XFILLER_52_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08428_ _08413_/A _08428_/B vssd1 vssd1 vccd1 vccd1 _08428_/X sky130_fd_sc_hd__and2b_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ _08359_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _08363_/A sky130_fd_sc_hd__xor2_1
XFILLER_149_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ _11368_/Y _11364_/C _11366_/Y _11367_/X vssd1 vssd1 vccd1 vccd1 _11371_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10321_ _10314_/B _10319_/B _10164_/X vssd1 vssd1 vccd1 vccd1 _10322_/B sky130_fd_sc_hd__o21a_1
XFILLER_109_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13040_ _13053_/C vssd1 vssd1 vccd1 vccd1 _13062_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10252_ _10340_/A vssd1 vssd1 vccd1 vccd1 _10338_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10183_ _10183_/A vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14991_ _14989_/Y _14985_/C _14987_/Y _14988_/X vssd1 vssd1 vccd1 vccd1 _14992_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_59_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16730_ _16730_/A _07835_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
X_13942_ _14092_/A vssd1 vssd1 vccd1 vccd1 _14063_/A sky130_fd_sc_hd__buf_2
XFILLER_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13873_ _13927_/A _13873_/B _13877_/B vssd1 vssd1 vccd1 vccd1 _16315_/D sky130_fd_sc_hd__nor3_1
XFILLER_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15612_ _15812_/CLK _15612_/D vssd1 vssd1 vccd1 vccd1 _15612_/Q sky130_fd_sc_hd__dfxtp_1
X_12824_ _12847_/A _12824_/B _12824_/C vssd1 vssd1 vccd1 vccd1 _12825_/A sky130_fd_sc_hd__and3_1
X_16592_ _16607_/CLK _16592_/D vssd1 vssd1 vccd1 vccd1 _16592_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15543_ _16551_/CLK _15543_/D vssd1 vssd1 vccd1 vccd1 _15543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _12755_/A vssd1 vssd1 vccd1 vccd1 _16157_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _16009_/Q _11878_/B _11706_/C vssd1 vssd1 vccd1 vccd1 _11706_/Y sky130_fd_sc_hd__nand3_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _16570_/CLK _15474_/D vssd1 vssd1 vccd1 vccd1 _15474_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12686_/A vssd1 vssd1 vccd1 vccd1 _12911_/B sky130_fd_sc_hd__buf_2
X_14425_ _14425_/A vssd1 vssd1 vccd1 vccd1 _16394_/D sky130_fd_sc_hd__clkbuf_1
X_11637_ _16001_/Q _11648_/C _11471_/X vssd1 vssd1 vccd1 vccd1 _11637_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14356_ _16386_/Q _14358_/C _14132_/X vssd1 vssd1 vccd1 vccd1 _14356_/Y sky130_fd_sc_hd__a21oi_1
X_11568_ _11569_/B _11569_/C _11567_/X vssd1 vssd1 vccd1 vccd1 _11570_/B sky130_fd_sc_hd__o21ai_1
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ _13304_/Y _13313_/A _13306_/Y _13302_/C vssd1 vssd1 vccd1 vccd1 _13309_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10519_ _10519_/A _10519_/B vssd1 vssd1 vccd1 vccd1 _10520_/B sky130_fd_sc_hd__nor2_1
X_14287_ _14851_/A vssd1 vssd1 vccd1 vccd1 _14287_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11499_ _15981_/Q _11500_/C _11441_/X vssd1 vssd1 vccd1 vccd1 _11501_/A sky130_fd_sc_hd__a21oi_1
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16026_ _16118_/CLK _16026_/D vssd1 vssd1 vccd1 vccd1 _16026_/Q sky130_fd_sc_hd__dfxtp_1
X_13238_ _13246_/A _13238_/B _13238_/C vssd1 vssd1 vccd1 vccd1 _13239_/A sky130_fd_sc_hd__and3_1
XFILLER_124_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13169_ _14015_/A vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09400_ _09400_/A vssd1 vssd1 vccd1 vccd1 _09497_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09331_ _09325_/C _09326_/C _09328_/Y _09335_/A vssd1 vssd1 vccd1 vccd1 _09335_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_80_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _09367_/A _09262_/B _09262_/C vssd1 vssd1 vccd1 vccd1 _09263_/A sky130_fd_sc_hd__and3_1
X_08213_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08225_/A sky130_fd_sc_hd__xor2_2
XFILLER_119_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09193_ _09193_/A _09193_/B vssd1 vssd1 vccd1 vccd1 _09195_/A sky130_fd_sc_hd__or2_1
XFILLER_119_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08144_ _08144_/A _08318_/A vssd1 vssd1 vccd1 vccd1 _08319_/A sky130_fd_sc_hd__xor2_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08075_ _08075_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08076_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08977_ _15531_/Q _08978_/C _08805_/X vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__a21o_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07928_ _07928_/A _07928_/B vssd1 vssd1 vccd1 vccd1 _07929_/B sky130_fd_sc_hd__nand2_1
X_07859_ _15552_/Q vssd1 vssd1 vccd1 vccd1 _08113_/A sky130_fd_sc_hd__inv_2
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ _10867_/Y _10880_/A _10869_/Y _10864_/C vssd1 vssd1 vccd1 vccd1 _10872_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09749_/A vssd1 vssd1 vccd1 vccd1 _09529_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12540_ _12540_/A _12540_/B _12540_/C vssd1 vssd1 vccd1 vccd1 _12541_/C sky130_fd_sc_hd__nand3_1
XFILLER_40_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _12505_/A _12471_/B _12471_/C vssd1 vssd1 vccd1 vccd1 _12472_/A sky130_fd_sc_hd__and3_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14210_ _14210_/A vssd1 vssd1 vccd1 vccd1 _14437_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11422_ _11420_/Y _11415_/C _11417_/Y _11419_/X vssd1 vssd1 vccd1 vccd1 _11423_/C
+ sky130_fd_sc_hd__a211o_1
X_15190_ _15184_/C _15185_/C _15187_/Y _15188_/X vssd1 vssd1 vccd1 vccd1 _15191_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14141_ _16355_/Q _14193_/B _14148_/C vssd1 vssd1 vccd1 vccd1 _14141_/X sky130_fd_sc_hd__and3_1
X_11353_ _15961_/Q _11353_/B _11353_/C vssd1 vssd1 vccd1 vccd1 _11353_/X sky130_fd_sc_hd__and3_1
XFILLER_4_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _10338_/A _10304_/B _10304_/C vssd1 vssd1 vccd1 vccd1 _10305_/A sky130_fd_sc_hd__and3_1
X_14072_ _16345_/Q _14179_/B _14072_/C vssd1 vssd1 vccd1 vccd1 _14072_/X sky130_fd_sc_hd__and3_1
X_11284_ _11452_/A _11284_/B _11284_/C vssd1 vssd1 vccd1 vccd1 _11285_/C sky130_fd_sc_hd__or3_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13023_ _16195_/Q _13194_/B _13028_/C vssd1 vssd1 vccd1 vccd1 _13023_/Y sky130_fd_sc_hd__nand3_1
X_10235_ _15780_/Q _10483_/B _10235_/C vssd1 vssd1 vccd1 vccd1 _10240_/A sky130_fd_sc_hd__and3_1
XFILLER_121_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10166_ _10322_/A _10166_/B vssd1 vssd1 vccd1 vccd1 _10166_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10097_ _10097_/A vssd1 vssd1 vccd1 vccd1 _15754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14974_ _16482_/Q _15027_/B _14974_/C vssd1 vssd1 vccd1 vccd1 _14974_/X sky130_fd_sc_hd__and3_1
XFILLER_75_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16713_ _16713_/A _07816_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_47_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13925_ _13920_/Y _13931_/A _13924_/Y _13918_/C vssd1 vssd1 vccd1 vccd1 _13927_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13856_ _16313_/Q _13856_/B _13856_/C vssd1 vssd1 vccd1 vccd1 _13856_/Y sky130_fd_sc_hd__nand3_1
XFILLER_34_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12807_ _12808_/B _12808_/C _12699_/X vssd1 vssd1 vccd1 vccd1 _12809_/B sky130_fd_sc_hd__o21ai_1
X_13787_ _16304_/Q _14010_/B _13793_/C vssd1 vssd1 vccd1 vccd1 _13789_/C sky130_fd_sc_hd__nand3_1
X_16575_ _16595_/CLK _16575_/D vssd1 vssd1 vccd1 vccd1 _16575_/Q sky130_fd_sc_hd__dfxtp_1
X_10999_ _11850_/A vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__buf_2
X_15526_ _15791_/CLK _15526_/D vssd1 vssd1 vccd1 vccd1 _15526_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _16156_/Q _12745_/C _12567_/X vssd1 vssd1 vccd1 vccd1 _12738_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15457_ _16551_/CLK _15457_/D vssd1 vssd1 vccd1 vccd1 _15457_/Q sky130_fd_sc_hd__dfxtp_2
X_12669_ _16146_/Q _12776_/B _12670_/C vssd1 vssd1 vccd1 vccd1 _12669_/X sky130_fd_sc_hd__and3_1
X_14408_ _14402_/C _14403_/C _14405_/Y _14406_/X vssd1 vssd1 vccd1 vccd1 _14409_/C
+ sky130_fd_sc_hd__a211o_1
X_15388_ _16013_/Q _16012_/Q _16011_/Q _15385_/X vssd1 vssd1 vccd1 vccd1 _16572_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14339_ _14906_/A vssd1 vssd1 vccd1 vccd1 _14339_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08900_ _08900_/A vssd1 vssd1 vccd1 vccd1 _15509_/D sky130_fd_sc_hd__clkbuf_1
X_16009_ _16554_/Q _16009_/D vssd1 vssd1 vccd1 vccd1 _16009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09880_/A _09880_/B vssd1 vssd1 vccd1 vccd1 _09880_/X sky130_fd_sc_hd__or2_1
XFILLER_98_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08831_/A _08836_/C vssd1 vssd1 vccd1 vccd1 _08835_/A sky130_fd_sc_hd__and2_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08846_/A _08762_/B _08768_/A vssd1 vssd1 vccd1 vccd1 _15481_/D sky130_fd_sc_hd__nor3_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08693_ _08693_/A _08693_/B vssd1 vssd1 vccd1 vccd1 _08694_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09314_ _09756_/A vssd1 vssd1 vccd1 vccd1 _09314_/X sky130_fd_sc_hd__buf_2
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09245_ _09125_/X _09243_/A _08667_/A vssd1 vssd1 vccd1 vccd1 _09246_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09176_ _09812_/A vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08127_ _14960_/A _07873_/B _07872_/B vssd1 vssd1 vccd1 vccd1 _08129_/C sky130_fd_sc_hd__o21a_1
XFILLER_107_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08058_ _08058_/A _08058_/B vssd1 vssd1 vccd1 vccd1 _08059_/B sky130_fd_sc_hd__nand2_2
XFILLER_134_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10020_ _09851_/X _10017_/B _10019_/Y vssd1 vssd1 vccd1 vccd1 _15739_/D sky130_fd_sc_hd__o21a_1
XFILLER_102_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11971_ _16048_/Q _11979_/C _11748_/X vssd1 vssd1 vccd1 vccd1 _11974_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13710_ _13710_/A _13717_/B vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__or2_1
X_10922_ _15898_/Q _10922_/B _10928_/C vssd1 vssd1 vccd1 vccd1 _10922_/Y sky130_fd_sc_hd__nand3_1
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14690_ _14688_/Y _14689_/X _14685_/C _14686_/C vssd1 vssd1 vccd1 vccd1 _14692_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13641_ _13637_/Y _13647_/A _13640_/Y _13635_/C vssd1 vssd1 vccd1 vccd1 _13643_/B
+ sky130_fd_sc_hd__o211a_1
X_10853_ _10849_/Y _10851_/X _10852_/Y _10847_/C vssd1 vssd1 vccd1 vccd1 _10855_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16389_/CLK _16360_/D vssd1 vssd1 vccd1 vccd1 _16360_/Q sky130_fd_sc_hd__dfxtp_1
X_13572_ _16274_/Q _13623_/B _13573_/C vssd1 vssd1 vccd1 vccd1 _13572_/X sky130_fd_sc_hd__and3_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _10777_/C _10778_/C _10781_/Y _10782_/X vssd1 vssd1 vccd1 vccd1 _10785_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15311_ _15311_/A _15311_/B vssd1 vssd1 vccd1 vccd1 _15312_/B sky130_fd_sc_hd__nand2_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _13371_/A vssd1 vssd1 vccd1 vccd1 _12751_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16291_ _16346_/CLK _16291_/D vssd1 vssd1 vccd1 vccd1 _16291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _15240_/Y _15241_/X _15237_/C _15238_/C vssd1 vssd1 vccd1 vccd1 _15244_/B
+ sky130_fd_sc_hd__o211ai_1
X_12454_ _12454_/A vssd1 vssd1 vccd1 vccd1 _16114_/D sky130_fd_sc_hd__clkbuf_1
X_11405_ _15968_/Q _11465_/B _11412_/C vssd1 vssd1 vccd1 vccd1 _11407_/C sky130_fd_sc_hd__nand3_1
X_15173_ _16504_/Q _16503_/Q _16502_/Q _15172_/X vssd1 vssd1 vccd1 vccd1 _16514_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_126_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ _16106_/Q _12387_/C _12157_/X vssd1 vssd1 vccd1 vccd1 _12385_/Y sky130_fd_sc_hd__a21oi_1
X_14124_ _14145_/A _14124_/B _14124_/C vssd1 vssd1 vccd1 vccd1 _14125_/A sky130_fd_sc_hd__and3_1
X_11336_ _11452_/A _11336_/B _11336_/C vssd1 vssd1 vccd1 vccd1 _11337_/C sky130_fd_sc_hd__or3_1
XFILLER_113_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14055_ _14055_/A vssd1 vssd1 vccd1 vccd1 _16341_/D sky130_fd_sc_hd__clkbuf_1
X_11267_ _15948_/Q _11275_/C _11150_/X vssd1 vssd1 vccd1 vccd1 _11267_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13006_ _13006_/A vssd1 vssd1 vccd1 vccd1 _13006_/X sky130_fd_sc_hd__buf_2
X_10218_ _10271_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10218_/X sky130_fd_sc_hd__or2_1
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11198_ _11195_/Y _11196_/X _11197_/Y _11193_/C vssd1 vssd1 vccd1 vccd1 _11200_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_67_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10149_ _13183_/A vssd1 vssd1 vccd1 vccd1 _12968_/A sky130_fd_sc_hd__buf_6
XFILLER_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14957_ _14992_/A _14957_/B _14957_/C vssd1 vssd1 vccd1 vccd1 _14958_/A sky130_fd_sc_hd__and3_1
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13908_ _16321_/Q _14135_/B _13908_/C vssd1 vssd1 vccd1 vccd1 _13908_/Y sky130_fd_sc_hd__nand3_1
X_14888_ _14888_/A _14896_/B vssd1 vssd1 vccd1 vccd1 _14890_/A sky130_fd_sc_hd__or2_1
XFILLER_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13839_ _16311_/Q _13948_/B _13848_/C vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__and3_1
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16558_ _16595_/CLK _16558_/D vssd1 vssd1 vccd1 vccd1 _16558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15509_ _15791_/CLK _15509_/D vssd1 vssd1 vccd1 vccd1 _15509_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_148_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16489_ _16607_/CLK _16489_/D vssd1 vssd1 vccd1 vccd1 _16489_/Q sky130_fd_sc_hd__dfxtp_1
X_09030_ _09030_/A _09030_/B vssd1 vssd1 vccd1 vccd1 _09031_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09932_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09863_ _15709_/Q _09884_/C _09714_/X vssd1 vssd1 vccd1 vccd1 _09865_/B sky130_fd_sc_hd__a21oi_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08814_ _08812_/Y _08824_/A _08809_/C _08810_/C vssd1 vssd1 vccd1 vccd1 _08816_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09617_/X _09706_/X _09788_/B _09707_/X vssd1 vssd1 vccd1 vccd1 _09795_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08745_ _08745_/A _08745_/B vssd1 vssd1 vccd1 vccd1 _15477_/D sky130_fd_sc_hd__nor2_1
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _08730_/A _08676_/B _08680_/A vssd1 vssd1 vccd1 vccd1 _15463_/D sky130_fd_sc_hd__nor3_1
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ _09222_/C _09223_/C _09225_/Y _09233_/A vssd1 vssd1 vccd1 vccd1 _09233_/B
+ sky130_fd_sc_hd__a211oi_1
X_09159_ _09076_/X _09151_/B _09154_/B _09158_/Y vssd1 vssd1 vccd1 vccd1 _15566_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_107_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12170_ _12170_/A _12170_/B _12170_/C vssd1 vssd1 vccd1 vccd1 _12171_/A sky130_fd_sc_hd__and3_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11121_ _15928_/Q _11183_/B _11128_/C vssd1 vssd1 vccd1 vccd1 _11123_/C sky130_fd_sc_hd__nand3_1
XFILLER_122_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11052_ _11053_/B _11053_/C _10999_/X vssd1 vssd1 vccd1 vccd1 _11054_/B sky130_fd_sc_hd__o21ai_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10003_ _15739_/Q _10003_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10005_/B sky130_fd_sc_hd__and3_1
XFILLER_1_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15860_ _16595_/CLK _15860_/D vssd1 vssd1 vccd1 vccd1 _15860_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14811_ _14819_/A _14811_/B _14811_/C vssd1 vssd1 vccd1 vccd1 _14812_/A sky130_fd_sc_hd__and3_1
X_15791_ _15791_/CLK _15791_/D vssd1 vssd1 vccd1 vccd1 _15791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11954_ _11954_/A _11954_/B vssd1 vssd1 vccd1 vccd1 _11960_/C sky130_fd_sc_hd__nor2_1
X_14742_ _16446_/Q _14742_/B _14742_/C vssd1 vssd1 vccd1 vccd1 _14742_/X sky130_fd_sc_hd__and3_1
XFILLER_72_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10905_ _13060_/A vssd1 vssd1 vccd1 vccd1 _10905_/X sky130_fd_sc_hd__buf_2
XFILLER_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14673_ _14673_/A vssd1 vssd1 vccd1 vccd1 _16432_/D sky130_fd_sc_hd__clkbuf_1
X_11885_ _16034_/Q _12053_/B _11891_/C vssd1 vssd1 vccd1 vccd1 _11885_/Y sky130_fd_sc_hd__nand3_1
XFILLER_83_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16412_ input11/X _16412_/D vssd1 vssd1 vccd1 vccd1 _16412_/Q sky130_fd_sc_hd__dfxtp_1
X_13624_ _14186_/A vssd1 vssd1 vccd1 vccd1 _13856_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10836_ _15888_/Q _10900_/B _10844_/C vssd1 vssd1 vccd1 vccd1 _10838_/C sky130_fd_sc_hd__nand3_1
Xrepeater22 _15812_/CLK vssd1 vssd1 vccd1 vccd1 _16595_/CLK sky130_fd_sc_hd__buf_12
X_13555_ _16271_/Q _13592_/C _13495_/X vssd1 vssd1 vccd1 vccd1 _13557_/B sky130_fd_sc_hd__a21oi_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16343_ _16389_/CLK _16343_/D vssd1 vssd1 vccd1 vccd1 _16343_/Q sky130_fd_sc_hd__dfxtp_1
X_10767_ _10767_/A vssd1 vssd1 vccd1 vccd1 _10782_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12506_ _12506_/A vssd1 vssd1 vccd1 vccd1 _16122_/D sky130_fd_sc_hd__clkbuf_1
X_16274_ _16533_/Q _16274_/D vssd1 vssd1 vccd1 vccd1 _16274_/Q sky130_fd_sc_hd__dfxtp_1
X_13486_ _13488_/B _13488_/C _13264_/X vssd1 vssd1 vccd1 vccd1 _13489_/B sky130_fd_sc_hd__o21ai_1
X_10698_ _11266_/A vssd1 vssd1 vccd1 vccd1 _10809_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15225_ _15225_/A vssd1 vssd1 vccd1 vccd1 _16522_/D sky130_fd_sc_hd__clkbuf_1
X_12437_ _12431_/C _12432_/C _12434_/Y _12435_/X vssd1 vssd1 vccd1 vccd1 _12438_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15156_ _16511_/Q _15156_/B _15161_/C vssd1 vssd1 vccd1 vccd1 _15156_/Y sky130_fd_sc_hd__nand3_1
X_12368_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__buf_2
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _14160_/A vssd1 vssd1 vccd1 vccd1 _14145_/A sky130_fd_sc_hd__clkbuf_2
X_11319_ _11319_/A _11319_/B _11319_/C vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__and3_1
X_15087_ _15087_/A vssd1 vssd1 vccd1 vccd1 _16499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12299_ _12299_/A _12299_/B vssd1 vssd1 vccd1 vccd1 _12304_/C sky130_fd_sc_hd__nor2_1
XFILLER_141_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14038_ _16340_/Q _14148_/B _14038_/C vssd1 vssd1 vccd1 vccd1 _14046_/A sky130_fd_sc_hd__and3_1
XFILLER_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15989_ _16005_/CLK _15989_/D vssd1 vssd1 vccd1 vccd1 _15989_/Q sky130_fd_sc_hd__dfxtp_1
X_08530_ _15312_/A _08530_/B vssd1 vssd1 vccd1 vccd1 _08530_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08461_ _08461_/A _08461_/B vssd1 vssd1 vccd1 vccd1 _08462_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08392_ _08393_/A _08393_/B vssd1 vssd1 vccd1 vccd1 _08394_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ _09054_/A _09013_/B _09018_/A vssd1 vssd1 vccd1 vccd1 _15535_/D sky130_fd_sc_hd__nor3_1
XFILLER_136_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09915_ _09913_/Y _09920_/A _09910_/C _09911_/C vssd1 vssd1 vccd1 vccd1 _09917_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09846_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__or2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09777_/X sky130_fd_sc_hd__or2_1
XFILLER_37_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08728_ _08726_/Y _08734_/A _08723_/C _08724_/C vssd1 vssd1 vccd1 vccd1 _08730_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _15274_/A vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__buf_2
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11670_/A _11670_/B vssd1 vssd1 vccd1 vccd1 _11673_/B sky130_fd_sc_hd__nor2_1
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10621_ _10469_/X _10613_/B _10616_/B _10620_/Y vssd1 vssd1 vccd1 vccd1 _15847_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13340_ _13340_/A vssd1 vssd1 vccd1 vccd1 _16240_/D sky130_fd_sc_hd__clkbuf_1
X_10552_ _15837_/Q _10691_/B _10559_/C vssd1 vssd1 vccd1 vccd1 _10552_/X sky130_fd_sc_hd__and3_1
XFILLER_128_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13271_ _13292_/C vssd1 vssd1 vccd1 vccd1 _13305_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10483_ _15825_/Q _10483_/B _10483_/C vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__and3_1
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15010_ _15045_/A _15010_/B _15010_/C vssd1 vssd1 vccd1 vccd1 _15011_/A sky130_fd_sc_hd__and3_1
X_12222_ _12222_/A _12222_/B _12222_/C vssd1 vssd1 vccd1 vccd1 _12223_/A sky130_fd_sc_hd__and3_1
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _12151_/Y _12152_/X _12148_/C _12149_/C vssd1 vssd1 vccd1 vccd1 _12155_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _11332_/A _11109_/C vssd1 vssd1 vccd1 vccd1 _11104_/X sky130_fd_sc_hd__or2_1
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12084_ _12084_/A _12084_/B _12089_/A vssd1 vssd1 vccd1 vccd1 _16062_/D sky130_fd_sc_hd__nor3_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11035_ _11033_/Y _11029_/C _11031_/Y _11032_/X vssd1 vssd1 vccd1 vccd1 _11036_/C
+ sky130_fd_sc_hd__a211o_1
X_15912_ _16553_/Q _15912_/D vssd1 vssd1 vccd1 vccd1 _15912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15843_ _16595_/CLK _15843_/D vssd1 vssd1 vccd1 vccd1 _15843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15774_ _15812_/CLK _15774_/D vssd1 vssd1 vccd1 vccd1 _15774_/Q sky130_fd_sc_hd__dfxtp_1
X_12986_ _12986_/A vssd1 vssd1 vccd1 vccd1 _16189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14725_ _14760_/A _14725_/B _14725_/C vssd1 vssd1 vccd1 vccd1 _14726_/A sky130_fd_sc_hd__and3_1
XFILLER_18_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11937_ _16042_/Q _12053_/B _11944_/C vssd1 vssd1 vccd1 vccd1 _11937_/Y sky130_fd_sc_hd__nand3_1
XFILLER_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11868_ _16033_/Q _11878_/C _11755_/X vssd1 vssd1 vccd1 vccd1 _11868_/Y sky130_fd_sc_hd__a21oi_1
X_14656_ _14941_/A vssd1 vssd1 vccd1 vccd1 _14882_/B sky130_fd_sc_hd__clkbuf_2
X_13607_ _16279_/Q _13645_/C _13495_/X vssd1 vssd1 vccd1 vccd1 _13609_/B sky130_fd_sc_hd__a21oi_1
X_10819_ _13652_/A vssd1 vssd1 vccd1 vccd1 _11957_/A sky130_fd_sc_hd__clkbuf_4
X_11799_ _11814_/C vssd1 vssd1 vccd1 vccd1 _11821_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14587_ _14587_/A vssd1 vssd1 vccd1 vccd1 _16419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16326_ _16346_/CLK _16326_/D vssd1 vssd1 vccd1 vccd1 _16326_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13538_ _16269_/Q _13645_/B _13538_/C vssd1 vssd1 vccd1 vccd1 _13548_/B sky130_fd_sc_hd__and3_1
XFILLER_145_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13469_ _13467_/Y _13462_/C _13465_/Y _13466_/X vssd1 vssd1 vccd1 vccd1 _13470_/C
+ sky130_fd_sc_hd__a211o_1
X_16257_ _16261_/CLK _16257_/D vssd1 vssd1 vccd1 vccd1 _16257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15208_ _16521_/Q _15215_/C _08747_/A vssd1 vssd1 vccd1 vccd1 _15208_/Y sky130_fd_sc_hd__a21oi_1
X_16188_ _16555_/Q _16188_/D vssd1 vssd1 vccd1 vccd1 _16188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15139_ _15139_/A vssd1 vssd1 vccd1 vccd1 _16508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07961_ _16581_/Q _16579_/Q vssd1 vssd1 vccd1 vccd1 _07963_/A sky130_fd_sc_hd__or2_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09700_ _09931_/A _09700_/B vssd1 vssd1 vccd1 vccd1 _09701_/B sky130_fd_sc_hd__and2_1
X_07892_ _07892_/A _07892_/B vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__xor2_4
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09631_ _09632_/B _09632_/C _09632_/A vssd1 vssd1 vccd1 vccd1 _09633_/B sky130_fd_sc_hd__a21o_1
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09562_ _15650_/Q _09561_/C _09383_/X vssd1 vssd1 vccd1 vccd1 _09563_/B sky130_fd_sc_hd__a21o_1
XFILLER_71_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08513_ _08472_/A _08472_/B _08512_/Y vssd1 vssd1 vccd1 vccd1 _08535_/B sky130_fd_sc_hd__a21oi_4
X_09493_ _09943_/A vssd1 vssd1 vccd1 vccd1 _09493_/X sky130_fd_sc_hd__buf_2
XFILLER_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08444_ _08444_/A _08444_/B vssd1 vssd1 vccd1 vccd1 _08445_/B sky130_fd_sc_hd__xnor2_2
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08375_ _08220_/A _08220_/B _08374_/Y vssd1 vssd1 vccd1 vccd1 _08377_/C sky130_fd_sc_hd__a21oi_2
XFILLER_149_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09829_ _09822_/Y _09826_/X _09828_/Y _09819_/C vssd1 vssd1 vccd1 vccd1 _09831_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _12840_/A vssd1 vssd1 vccd1 vccd1 _16169_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12769_/Y _12770_/X _12766_/C _12767_/C vssd1 vssd1 vccd1 vccd1 _12773_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _16011_/Q _11780_/B _11729_/C vssd1 vssd1 vccd1 vccd1 _11722_/Y sky130_fd_sc_hd__nand3_1
XFILLER_64_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14510_ _14511_/B _14511_/C _14511_/A vssd1 vssd1 vccd1 vccd1 _14512_/B sky130_fd_sc_hd__a21o_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _16570_/CLK _15490_/D vssd1 vssd1 vccd1 vccd1 _15490_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11653_ _16003_/Q _11662_/C _11485_/X vssd1 vssd1 vccd1 vccd1 _11653_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _14555_/A _14441_/B _14441_/C vssd1 vssd1 vccd1 vccd1 _14442_/C sky130_fd_sc_hd__or3_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10604_ _10604_/A vssd1 vssd1 vccd1 vccd1 _15844_/D sky130_fd_sc_hd__clkbuf_1
X_14372_ _16388_/Q _14380_/C _14258_/X vssd1 vssd1 vccd1 vccd1 _14372_/Y sky130_fd_sc_hd__a21oi_1
X_11584_ _11584_/A vssd1 vssd1 vccd1 vccd1 _15991_/D sky130_fd_sc_hd__clkbuf_1
X_13323_ _13336_/C vssd1 vssd1 vccd1 vccd1 _13344_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _16118_/CLK _16111_/D vssd1 vssd1 vccd1 vccd1 _16111_/Q sky130_fd_sc_hd__dfxtp_1
X_10535_ _10833_/B vssd1 vssd1 vccd1 vccd1 _10726_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16042_ _16118_/CLK _16042_/D vssd1 vssd1 vccd1 vccd1 _16042_/Q sky130_fd_sc_hd__dfxtp_1
X_13254_ _13252_/Y _13246_/C _13249_/Y _13259_/A vssd1 vssd1 vccd1 vccd1 _13259_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ _10466_/A _10466_/B vssd1 vssd1 vccd1 vccd1 _10467_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12205_ _12203_/Y _12204_/X _12200_/C _12201_/C vssd1 vssd1 vccd1 vccd1 _12207_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _16219_/Q _13193_/C _13184_/X vssd1 vssd1 vccd1 vccd1 _13185_/Y sky130_fd_sc_hd__a21oi_1
X_10397_ _10394_/Y _10395_/X _10396_/Y _10391_/C vssd1 vssd1 vccd1 vccd1 _10399_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12136_ _12170_/A _12136_/B _12136_/C vssd1 vssd1 vccd1 vccd1 _12137_/A sky130_fd_sc_hd__and3_1
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12067_ _12067_/A _12067_/B vssd1 vssd1 vccd1 vccd1 _12068_/B sky130_fd_sc_hd__nor2_1
X_11018_ _15913_/Q _11070_/B _11018_/C vssd1 vssd1 vccd1 vccd1 _11018_/X sky130_fd_sc_hd__and3_1
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15826_ _16570_/CLK _15826_/D vssd1 vssd1 vccd1 vccd1 _15826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15757_ _15812_/CLK _15757_/D vssd1 vssd1 vccd1 vccd1 _15757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12969_ _14095_/A vssd1 vssd1 vccd1 vccd1 _13194_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14708_ _14708_/A vssd1 vssd1 vccd1 vccd1 _16438_/D sky130_fd_sc_hd__clkbuf_1
X_15688_ _15791_/CLK _15688_/D vssd1 vssd1 vccd1 vccd1 _15688_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ _16429_/Q _14748_/B _14640_/C vssd1 vssd1 vccd1 vccd1 _14639_/X sky130_fd_sc_hd__and3_1
XFILLER_21_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08160_ _08160_/A _08331_/A vssd1 vssd1 vccd1 vccd1 _08176_/A sky130_fd_sc_hd__xnor2_1
X_16309_ _16346_/CLK _16309_/D vssd1 vssd1 vccd1 vccd1 _16309_/Q sky130_fd_sc_hd__dfxtp_1
X_08091_ _16564_/Q _08276_/B vssd1 vssd1 vccd1 vccd1 _08092_/B sky130_fd_sc_hd__xnor2_1
XFILLER_119_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08993_ _08993_/A _08993_/B vssd1 vssd1 vccd1 vccd1 _08994_/B sky130_fd_sc_hd__nor2_1
XFILLER_141_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07944_ _11798_/A _07944_/B vssd1 vssd1 vccd1 vccd1 _07945_/B sky130_fd_sc_hd__xnor2_2
XFILLER_56_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07875_ _12928_/A _07876_/B vssd1 vssd1 vccd1 vccd1 _07877_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09614_ _09529_/X _09611_/B _09613_/Y vssd1 vssd1 vccd1 vccd1 _15658_/D sky130_fd_sc_hd__o21a_1
XFILLER_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _09546_/B _09546_/C _09546_/A vssd1 vssd1 vccd1 vccd1 _09547_/B sky130_fd_sc_hd__a21o_1
XFILLER_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09476_ _09471_/Y _09474_/X _09475_/Y vssd1 vssd1 vccd1 vccd1 _15629_/D sky130_fd_sc_hd__o21a_1
X_08427_ _15221_/A vssd1 vssd1 vccd1 vccd1 _15304_/A sky130_fd_sc_hd__clkbuf_4
X_08358_ _08213_/A _08213_/B _08356_/X _08357_/Y vssd1 vssd1 vccd1 vccd1 _08359_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08289_ _08098_/A _08098_/B _08288_/Y vssd1 vssd1 vccd1 vccd1 _08408_/B sky130_fd_sc_hd__o21a_1
XFILLER_137_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10320_ _10318_/A _10318_/B _10319_/X vssd1 vssd1 vccd1 vccd1 _15792_/D sky130_fd_sc_hd__a21oi_1
XFILLER_124_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _10251_/A vssd1 vssd1 vccd1 vccd1 _15780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _15772_/Q _10190_/C _10181_/X vssd1 vssd1 vccd1 vccd1 _10186_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14990_ _14987_/Y _14988_/X _14989_/Y _14985_/C vssd1 vssd1 vccd1 vccd1 _14992_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13941_ _13941_/A vssd1 vssd1 vccd1 vccd1 _16325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13872_ _13870_/Y _13866_/C _13868_/Y _13877_/A vssd1 vssd1 vccd1 vccd1 _13877_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ _15812_/CLK _15611_/D vssd1 vssd1 vccd1 vccd1 _15611_/Q sky130_fd_sc_hd__dfxtp_1
X_12823_ _12823_/A _12823_/B _12823_/C vssd1 vssd1 vccd1 vccd1 _12824_/C sky130_fd_sc_hd__nand3_1
XFILLER_15_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16591_ _16607_/CLK _16591_/D vssd1 vssd1 vccd1 vccd1 _16591_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15542_ _16551_/CLK _15542_/D vssd1 vssd1 vccd1 vccd1 _15542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12788_/A _12754_/B _12754_/C vssd1 vssd1 vccd1 vccd1 _12755_/A sky130_fd_sc_hd__and3_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11705_ _16010_/Q _11928_/B _11706_/C vssd1 vssd1 vccd1 vccd1 _11705_/X sky130_fd_sc_hd__and3_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15473_ _16570_/CLK _15473_/D vssd1 vssd1 vccd1 vccd1 _15473_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _16148_/Q _12739_/B _12685_/C vssd1 vssd1 vccd1 vccd1 _12694_/A sky130_fd_sc_hd__and3_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ _11636_/A vssd1 vssd1 vccd1 vccd1 _15999_/D sky130_fd_sc_hd__clkbuf_1
X_14424_ _14424_/A _14424_/B _14424_/C vssd1 vssd1 vccd1 vccd1 _14425_/A sky130_fd_sc_hd__and3_1
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _11850_/A vssd1 vssd1 vccd1 vccd1 _11567_/X sky130_fd_sc_hd__clkbuf_2
X_14355_ _14355_/A vssd1 vssd1 vccd1 vccd1 _16384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10518_ _10518_/A _10518_/B vssd1 vssd1 vccd1 vccd1 _10520_/A sky130_fd_sc_hd__or2_1
X_13306_ _16235_/Q _13474_/B _13311_/C vssd1 vssd1 vccd1 vccd1 _13306_/Y sky130_fd_sc_hd__nand3_1
X_14286_ _14342_/A _14286_/B _14291_/A vssd1 vssd1 vccd1 vccd1 _16374_/D sky130_fd_sc_hd__nor3_1
X_11498_ _11520_/A _11498_/B _11502_/B vssd1 vssd1 vccd1 vccd1 _15979_/D sky130_fd_sc_hd__nor3_1
XFILLER_109_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16025_ _16118_/CLK _16025_/D vssd1 vssd1 vccd1 vccd1 _16025_/Q sky130_fd_sc_hd__dfxtp_1
X_13237_ _13235_/Y _13231_/C _13233_/Y _13234_/X vssd1 vssd1 vccd1 vccd1 _13238_/C
+ sky130_fd_sc_hd__a211o_1
X_10449_ _10445_/Y _10446_/X _10448_/Y _10443_/C vssd1 vssd1 vccd1 vccd1 _10451_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13168_ _13168_/A vssd1 vssd1 vccd1 vccd1 _16215_/D sky130_fd_sc_hd__clkbuf_1
X_12119_ _12686_/A vssd1 vssd1 vccd1 vccd1 _12347_/B sky130_fd_sc_hd__clkbuf_2
X_13099_ _13120_/C vssd1 vssd1 vccd1 vccd1 _13135_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15809_ _16570_/CLK _15809_/D vssd1 vssd1 vccd1 vccd1 _15809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _09328_/Y _09335_/A _09325_/C _09326_/C vssd1 vssd1 vccd1 vccd1 _09332_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09261_ _09261_/A _09261_/B _09261_/C vssd1 vssd1 vccd1 vccd1 _09262_/C sky130_fd_sc_hd__nand3_1
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08212_ _08357_/B _08212_/B vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__nor2_1
X_09192_ _15578_/Q _09192_/B _09192_/C vssd1 vssd1 vccd1 vccd1 _09193_/B sky130_fd_sc_hd__and3_1
X_08143_ _08143_/A _08143_/B vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__xnor2_1
XFILLER_147_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08074_ _15579_/Q _15561_/Q vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__or2_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08976_ _09812_/A vssd1 vssd1 vccd1 vccd1 _09142_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07927_ _16598_/Q _16596_/Q vssd1 vssd1 vccd1 vccd1 _07928_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07858_ _15516_/Q vssd1 vssd1 vccd1 vccd1 _08302_/A sky130_fd_sc_hd__inv_2
XFILLER_29_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07789_ _07793_/A vssd1 vssd1 vccd1 vccd1 _07789_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09528_ _09524_/X _09526_/B _09527_/Y vssd1 vssd1 vccd1 vccd1 _15639_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ _09456_/Y _09467_/A _09453_/C _09454_/C vssd1 vssd1 vccd1 vccd1 _09461_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12470_ _12586_/A _12470_/B _12470_/C vssd1 vssd1 vccd1 vccd1 _12471_/C sky130_fd_sc_hd__or3_1
XFILLER_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11421_ _11417_/Y _11419_/X _11420_/Y _11415_/C vssd1 vssd1 vccd1 vccd1 _11423_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14140_ _16355_/Q _14148_/C _14029_/X vssd1 vssd1 vccd1 vccd1 _14140_/Y sky130_fd_sc_hd__a21oi_1
X_11352_ _15961_/Q _11361_/C _11188_/X vssd1 vssd1 vccd1 vccd1 _11352_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10303_ _10301_/Y _10297_/C _10299_/Y _10300_/X vssd1 vssd1 vccd1 vccd1 _10304_/C
+ sky130_fd_sc_hd__a211o_1
X_14071_ _16345_/Q _14079_/C _14015_/X vssd1 vssd1 vccd1 vccd1 _14071_/Y sky130_fd_sc_hd__a21oi_1
X_11283_ _11284_/B _11284_/C _11282_/X vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__o21ai_1
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13022_ _16196_/Q _13022_/B _13022_/C vssd1 vssd1 vccd1 vccd1 _13030_/A sky130_fd_sc_hd__and3_1
X_10234_ _10833_/B vssd1 vssd1 vccd1 vccd1 _10483_/B sky130_fd_sc_hd__clkbuf_2
X_10165_ _10159_/B _10162_/B _10164_/X vssd1 vssd1 vccd1 vccd1 _10166_/B sky130_fd_sc_hd__o21a_1
XFILLER_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10096_ _10145_/A _10096_/B _10096_/C vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__and3_1
X_14973_ _16482_/Q _14982_/C _14858_/X vssd1 vssd1 vccd1 vccd1 _14973_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16712_ _16712_/A _07815_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
X_13924_ _16323_/Q _14039_/B _13929_/C vssd1 vssd1 vccd1 vccd1 _13924_/Y sky130_fd_sc_hd__nand3_1
XFILLER_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855_ _16314_/Q _13906_/B _13856_/C vssd1 vssd1 vccd1 vccd1 _13855_/X sky130_fd_sc_hd__and3_1
XFILLER_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ _13034_/A vssd1 vssd1 vccd1 vccd1 _12847_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16574_ _16595_/CLK _16574_/D vssd1 vssd1 vccd1 vccd1 _16574_/Q sky130_fd_sc_hd__dfxtp_1
X_13786_ _13786_/A vssd1 vssd1 vccd1 vccd1 _14010_/B sky130_fd_sc_hd__buf_2
X_10998_ _11051_/A vssd1 vssd1 vccd1 vccd1 _11036_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15525_ _16551_/CLK _15525_/D vssd1 vssd1 vccd1 vccd1 _15525_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12737_/A vssd1 vssd1 vccd1 vccd1 _16154_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15456_ _16570_/CLK _15456_/D vssd1 vssd1 vccd1 vccd1 _15456_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_129_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ _16146_/Q _12670_/C _12440_/X vssd1 vssd1 vccd1 vccd1 _12668_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14407_ _14405_/Y _14406_/X _14402_/C _14403_/C vssd1 vssd1 vccd1 vccd1 _14409_/B
+ sky130_fd_sc_hd__o211ai_1
X_11619_ _11619_/A vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15387_ _16005_/Q _16004_/Q _16003_/Q _15385_/X vssd1 vssd1 vccd1 vccd1 _16571_/D
+ sky130_fd_sc_hd__o31a_1
X_12599_ _16136_/Q _12607_/C _12598_/X vssd1 vssd1 vccd1 vccd1 _12602_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14338_ _14373_/C vssd1 vssd1 vccd1 vccd1 _14380_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14269_ _14269_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _14271_/A sky130_fd_sc_hd__or2_1
X_16008_ _16554_/Q _16008_/D vssd1 vssd1 vccd1 vccd1 _16008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _08630_/X _08823_/B _08826_/B _08829_/Y vssd1 vssd1 vccd1 vccd1 _15494_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _15485_/Q _08845_/B _08766_/C vssd1 vssd1 vccd1 vccd1 _08768_/A sky130_fd_sc_hd__and3_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08692_ _10060_/A vssd1 vssd1 vccd1 vccd1 _08870_/A sky130_fd_sc_hd__buf_2
XFILLER_66_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09313_ _09313_/A _09313_/B vssd1 vssd1 vccd1 vccd1 _15596_/D sky130_fd_sc_hd__nor2_1
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09244_ _15358_/A _15358_/B _09244_/C vssd1 vssd1 vccd1 vccd1 _09246_/A sky130_fd_sc_hd__and3_1
XFILLER_22_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09175_ _09256_/A _09175_/B _09180_/A vssd1 vssd1 vccd1 vccd1 _15571_/D sky130_fd_sc_hd__nor3_1
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08126_ _11683_/A _07914_/B _07917_/A vssd1 vssd1 vccd1 vccd1 _08136_/A sky130_fd_sc_hd__o21ai_4
XFILLER_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08057_ _15687_/Q _15669_/Q vssd1 vssd1 vccd1 vccd1 _08058_/B sky130_fd_sc_hd__or2_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08959_ _08832_/X _08963_/C _08924_/X vssd1 vssd1 vccd1 vccd1 _08960_/B sky130_fd_sc_hd__o21ai_1
X_16665__70 vssd1 vssd1 vccd1 vccd1 _16665__70/HI _16741_/A sky130_fd_sc_hd__conb_1
XFILLER_69_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11970_ _12084_/A _11970_/B _11974_/A vssd1 vssd1 vccd1 vccd1 _16046_/D sky130_fd_sc_hd__nor3_1
XFILLER_56_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10921_ _15899_/Q _11084_/B _10928_/C vssd1 vssd1 vccd1 vccd1 _10921_/X sky130_fd_sc_hd__and3_1
XFILLER_112_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10852_ _15889_/Q _11026_/B _10852_/C vssd1 vssd1 vccd1 vccd1 _10852_/Y sky130_fd_sc_hd__nand3_1
X_13640_ _16283_/Q _13760_/B _13645_/C vssd1 vssd1 vccd1 vccd1 _13640_/Y sky130_fd_sc_hd__nand3_1
XFILLER_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10781_/Y _10782_/X _10777_/C _10778_/C vssd1 vssd1 vccd1 vccd1 _10785_/B
+ sky130_fd_sc_hd__o211ai_1
X_13571_ _16274_/Q _13573_/C _13570_/X vssd1 vssd1 vccd1 vccd1 _13571_/Y sky130_fd_sc_hd__a21oi_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _15301_/A _15303_/B _15300_/A vssd1 vssd1 vccd1 vccd1 _15311_/B sky130_fd_sc_hd__a21o_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12520_/A _12520_/B _12521_/X vssd1 vssd1 vccd1 vccd1 _16124_/D sky130_fd_sc_hd__a21oi_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16533_/Q _16290_/D vssd1 vssd1 vccd1 vccd1 _16290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _16527_/Q _15241_/B _15241_/C vssd1 vssd1 vccd1 vccd1 _15241_/X sky130_fd_sc_hd__and3_1
X_12453_ _12453_/A _12453_/B _12453_/C vssd1 vssd1 vccd1 vccd1 _12454_/A sky130_fd_sc_hd__and3_1
X_11404_ _15968_/Q _11412_/C _11181_/X vssd1 vssd1 vccd1 vccd1 _11407_/B sky130_fd_sc_hd__a21o_1
X_15172_ _15378_/A vssd1 vssd1 vccd1 vccd1 _15172_/X sky130_fd_sc_hd__buf_4
X_12384_ _12384_/A vssd1 vssd1 vccd1 vccd1 _16104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11335_ _11336_/B _11336_/C _11282_/X vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__o21ai_1
X_14123_ _14123_/A _14123_/B _14123_/C vssd1 vssd1 vccd1 vccd1 _14124_/C sky130_fd_sc_hd__nand3_1
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ _11266_/A vssd1 vssd1 vccd1 vccd1 _11379_/A sky130_fd_sc_hd__buf_2
X_14054_ _14090_/A _14054_/B _14054_/C vssd1 vssd1 vccd1 vccd1 _14055_/A sky130_fd_sc_hd__and3_1
XFILLER_140_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10217_ _10217_/A _10217_/B vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__nor2_1
X_13005_ _13005_/A vssd1 vssd1 vccd1 vccd1 _16192_/D sky130_fd_sc_hd__clkbuf_1
X_11197_ _15937_/Q _11309_/B _11197_/C vssd1 vssd1 vccd1 vccd1 _11197_/Y sky130_fd_sc_hd__nand3_1
XFILLER_95_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ input4/X vssd1 vssd1 vccd1 vccd1 _13183_/A sky130_fd_sc_hd__buf_2
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10079_ _15754_/Q _10288_/C _10086_/C vssd1 vssd1 vccd1 vccd1 _10081_/C sky130_fd_sc_hd__nand3_1
X_14956_ _15117_/A _14956_/B _14956_/C vssd1 vssd1 vccd1 vccd1 _14957_/C sky130_fd_sc_hd__or3_1
XFILLER_48_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13907_ _14186_/A vssd1 vssd1 vccd1 vccd1 _14135_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14887_ _16468_/Q _15055_/B _14887_/C vssd1 vssd1 vccd1 vccd1 _14896_/B sky130_fd_sc_hd__and3_1
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13838_ _16311_/Q _13875_/C _13781_/X vssd1 vssd1 vccd1 vccd1 _13840_/B sky130_fd_sc_hd__a21oi_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16557_ _16595_/CLK _16557_/D vssd1 vssd1 vccd1 vccd1 _16557_/Q sky130_fd_sc_hd__dfxtp_1
X_13769_ _13879_/A _13774_/C vssd1 vssd1 vccd1 vccd1 _13769_/X sky130_fd_sc_hd__or2_1
XFILLER_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15508_ _15791_/CLK _15508_/D vssd1 vssd1 vccd1 vccd1 _15508_/Q sky130_fd_sc_hd__dfxtp_2
X_16488_ _16607_/CLK _16488_/D vssd1 vssd1 vccd1 vccd1 _16488_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15439_ _16349_/Q _16348_/Q _16347_/Q _15434_/X vssd1 vssd1 vccd1 vccd1 _16614_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09931_ _09931_/A _09931_/B vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__and2_1
X_09862_ _09873_/C vssd1 vssd1 vccd1 vccd1 _09884_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _15496_/Q _08943_/B _08822_/C vssd1 vssd1 vccd1 vccd1 _08824_/A sky130_fd_sc_hd__and3_1
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09615_/X _09788_/B _09792_/X vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__a21oi_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08744_ _08644_/X _08752_/C _08708_/X vssd1 vssd1 vccd1 vccd1 _08745_/B sky130_fd_sc_hd__o21ai_1
XFILLER_73_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _15467_/Q _08845_/B _08678_/C vssd1 vssd1 vccd1 vccd1 _08680_/A sky130_fd_sc_hd__and3_1
XFILLER_26_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09227_ _09225_/Y _09233_/A _09222_/C _09223_/C vssd1 vssd1 vccd1 vccd1 _09229_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09158_ _10065_/A _09165_/C vssd1 vssd1 vccd1 vccd1 _09158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08109_ _15367_/B _08109_/B _08109_/C vssd1 vssd1 vccd1 vccd1 _15446_/D sky130_fd_sc_hd__nor3_1
X_09089_ _09087_/X _09086_/A _09088_/Y vssd1 vssd1 vccd1 vccd1 _15551_/D sky130_fd_sc_hd__o21a_1
XFILLER_107_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11120_ _15928_/Q _11128_/C _10898_/X vssd1 vssd1 vccd1 vccd1 _11123_/B sky130_fd_sc_hd__a21o_1
XFILLER_116_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _11051_/A vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10002_ _15739_/Q _10009_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _10005_/A sky130_fd_sc_hd__a21oi_1
XFILLER_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14810_ _14808_/Y _14803_/C _14805_/Y _14807_/X vssd1 vssd1 vccd1 vccd1 _14811_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15790_ _15791_/CLK _15790_/D vssd1 vssd1 vccd1 vccd1 _15790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14741_ _16446_/Q _14750_/C _14574_/X vssd1 vssd1 vccd1 vccd1 _14741_/Y sky130_fd_sc_hd__a21oi_1
X_11953_ _12801_/A vssd1 vssd1 vccd1 vccd1 _12183_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10904_ _10904_/A vssd1 vssd1 vccd1 vccd1 _15895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14672_ _14707_/A _14672_/B _14672_/C vssd1 vssd1 vccd1 vccd1 _14673_/A sky130_fd_sc_hd__and3_1
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11884_ _16035_/Q _11936_/B _11891_/C vssd1 vssd1 vccd1 vccd1 _11884_/X sky130_fd_sc_hd__and3_1
X_16411_ input11/X _16411_/D vssd1 vssd1 vccd1 vccd1 _16411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13623_ _16282_/Q _13623_/B _13625_/C vssd1 vssd1 vccd1 vccd1 _13623_/X sky130_fd_sc_hd__and3_1
X_10835_ _15888_/Q _10844_/C _15235_/B vssd1 vssd1 vccd1 vccd1 _10838_/B sky130_fd_sc_hd__a21o_1
Xrepeater12 _15365_/A vssd1 vssd1 vccd1 vccd1 _16005_/CLK sky130_fd_sc_hd__buf_12
Xrepeater23 input11/X vssd1 vssd1 vccd1 vccd1 _16607_/CLK sky130_fd_sc_hd__buf_12
X_16342_ _16389_/CLK _16342_/D vssd1 vssd1 vccd1 vccd1 _16342_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _13586_/C vssd1 vssd1 vccd1 vccd1 _13592_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_9_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10766_ _15866_/Q _15865_/Q _15864_/Q _10719_/X vssd1 vssd1 vccd1 vccd1 _15876_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_9_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ _12505_/A _12505_/B _12505_/C vssd1 vssd1 vccd1 vccd1 _12506_/A sky130_fd_sc_hd__and3_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16273_ _16533_/Q _16273_/D vssd1 vssd1 vccd1 vccd1 _16273_/Q sky130_fd_sc_hd__dfxtp_1
X_10697_ _10697_/A vssd1 vssd1 vccd1 vccd1 _11266_/A sky130_fd_sc_hd__buf_4
X_13485_ _13598_/A vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15224_ _15258_/A _15224_/B _15224_/C vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__and3_1
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12436_ _12434_/Y _12435_/X _12431_/C _12432_/C vssd1 vssd1 vccd1 vccd1 _12438_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15155_ _16512_/Q _15261_/B _15155_/C vssd1 vssd1 vccd1 vccd1 _15163_/A sky130_fd_sc_hd__and3_1
X_12367_ _12402_/C vssd1 vssd1 vccd1 vccd1 _12409_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_114_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14106_ _14104_/A _14104_/B _14105_/X vssd1 vssd1 vccd1 vccd1 _16348_/D sky130_fd_sc_hd__a21oi_1
X_11318_ _11316_/Y _11312_/C _11314_/Y _11315_/X vssd1 vssd1 vccd1 vccd1 _11319_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15086_ _15100_/A _15086_/B _15086_/C vssd1 vssd1 vccd1 vccd1 _15087_/A sky130_fd_sc_hd__and3_1
X_12298_ _12298_/A _12298_/B vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__nor2_1
XFILLER_141_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11249_ _11264_/A _11249_/B _11249_/C vssd1 vssd1 vccd1 vccd1 _11250_/A sky130_fd_sc_hd__and3_1
X_14037_ _16340_/Q _14044_/C _13979_/X vssd1 vssd1 vccd1 vccd1 _14037_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15988_ _16005_/CLK _15988_/D vssd1 vssd1 vccd1 vccd1 _15988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14939_ _16476_/Q _14947_/C _14821_/X vssd1 vssd1 vccd1 vccd1 _14939_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08460_ _08395_/A _08395_/B _08394_/A vssd1 vssd1 vccd1 vccd1 _08461_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16609_ input11/X _16609_/D vssd1 vssd1 vccd1 vccd1 _16609_/Q sky130_fd_sc_hd__dfxtp_1
X_08391_ _08275_/A _08275_/B _08274_/A vssd1 vssd1 vccd1 vccd1 _08393_/B sky130_fd_sc_hd__a21oi_1
XFILLER_149_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _15539_/Q _09053_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09018_/A sky130_fd_sc_hd__and3_1
XFILLER_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09914_ _15720_/Q _09914_/B _09914_/C vssd1 vssd1 vccd1 vccd1 _09920_/A sky130_fd_sc_hd__and3_1
XFILLER_120_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09845_ _15704_/Q _10313_/C _09845_/C vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__and3_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09776_ _09776_/A _09776_/B vssd1 vssd1 vccd1 vccd1 _09776_/Y sky130_fd_sc_hd__nor2_1
X_16635__40 vssd1 vssd1 vccd1 vccd1 _16635__40/HI _16701_/A sky130_fd_sc_hd__conb_1
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08727_ _15478_/Q _10743_/B _08732_/C vssd1 vssd1 vccd1 vccd1 _08734_/A sky130_fd_sc_hd__and3_1
XFILLER_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _14895_/A vssd1 vssd1 vccd1 vccd1 _15274_/A sky130_fd_sc_hd__buf_2
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08589_/A vssd1 vssd1 vccd1 vccd1 _08807_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10620_ _15353_/A _10620_/B vssd1 vssd1 vccd1 vccd1 _10620_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ _15837_/Q _10559_/C _10393_/X vssd1 vssd1 vccd1 vccd1 _10551_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13270_ _13283_/C vssd1 vssd1 vccd1 vccd1 _13292_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10482_ _15825_/Q _10517_/C _10426_/X vssd1 vssd1 vccd1 vccd1 _10484_/B sky130_fd_sc_hd__a21oi_1
XFILLER_148_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12221_ _12219_/Y _12215_/C _12217_/Y _12218_/X vssd1 vssd1 vccd1 vccd1 _12222_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ _16073_/Q _12204_/B _12152_/C vssd1 vssd1 vccd1 vccd1 _12152_/X sky130_fd_sc_hd__and3_1
XFILLER_118_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11103_ _11103_/A _11103_/B vssd1 vssd1 vccd1 vccd1 _11109_/C sky130_fd_sc_hd__nor2_1
XFILLER_123_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12083_ _16063_/Q _12252_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__and3_1
XFILLER_111_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11034_ _11031_/Y _11032_/X _11033_/Y _11029_/C vssd1 vssd1 vccd1 vccd1 _11036_/B
+ sky130_fd_sc_hd__o211ai_1
X_15911_ _15365_/A _15911_/D vssd1 vssd1 vccd1 vccd1 _15911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15842_ _16595_/CLK _15842_/D vssd1 vssd1 vccd1 vccd1 _15842_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15773_ _15791_/CLK _15773_/D vssd1 vssd1 vccd1 vccd1 _15773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ _13019_/A _12985_/B _12985_/C vssd1 vssd1 vccd1 vccd1 _12986_/A sky130_fd_sc_hd__and3_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14724_ _14839_/A _14724_/B _14724_/C vssd1 vssd1 vccd1 vccd1 _14725_/C sky130_fd_sc_hd__or3_1
X_11936_ _16043_/Q _11936_/B _11944_/C vssd1 vssd1 vccd1 vccd1 _11936_/X sky130_fd_sc_hd__and3_1
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14655_ _16431_/Q _14710_/B _14655_/C vssd1 vssd1 vccd1 vccd1 _14664_/A sky130_fd_sc_hd__and3_1
X_11867_ _11867_/A vssd1 vssd1 vccd1 vccd1 _16031_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _13639_/C vssd1 vssd1 vccd1 vccd1 _13645_/C sky130_fd_sc_hd__clkbuf_2
X_10818_ _10816_/A _10816_/B _10817_/X vssd1 vssd1 vccd1 vccd1 _15883_/D sky130_fd_sc_hd__a21oi_1
X_14586_ _14594_/A _14586_/B _14586_/C vssd1 vssd1 vccd1 vccd1 _14587_/A sky130_fd_sc_hd__and3_1
X_11798_ _11798_/A vssd1 vssd1 vccd1 vccd1 _11814_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16325_ _16346_/CLK _16325_/D vssd1 vssd1 vccd1 vccd1 _16325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13537_ _16269_/Q _13538_/C _13421_/X vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__a21oi_1
X_10749_ _15874_/Q _10929_/B _10749_/C vssd1 vssd1 vccd1 vccd1 _10757_/A sky130_fd_sc_hd__and3_1
XFILLER_146_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16256_ _16261_/CLK _16256_/D vssd1 vssd1 vccd1 vccd1 _16256_/Q sky130_fd_sc_hd__dfxtp_1
X_13468_ _13465_/Y _13466_/X _13467_/Y _13462_/C vssd1 vssd1 vccd1 vccd1 _13470_/B
+ sky130_fd_sc_hd__o211ai_1
X_15207_ _15207_/A vssd1 vssd1 vccd1 vccd1 _15333_/A sky130_fd_sc_hd__buf_4
X_12419_ _12453_/A _12419_/B _12419_/C vssd1 vssd1 vccd1 vccd1 _12420_/A sky130_fd_sc_hd__and3_1
X_16187_ _16555_/Q _16187_/D vssd1 vssd1 vccd1 vccd1 _16187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13399_ _13682_/A vssd1 vssd1 vccd1 vccd1 _13623_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15138_ _15152_/A _15138_/B _15138_/C vssd1 vssd1 vccd1 vccd1 _15139_/A sky130_fd_sc_hd__and3_1
XFILLER_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15069_ _15069_/A vssd1 vssd1 vccd1 vccd1 _15083_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_07960_ _16583_/Q vssd1 vssd1 vccd1 vccd1 _12307_/A sky130_fd_sc_hd__clkinv_2
XFILLER_141_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07891_ _16568_/Q _08124_/B vssd1 vssd1 vccd1 vccd1 _07892_/B sky130_fd_sc_hd__xnor2_4
X_09630_ _15665_/Q _09867_/B _09636_/C vssd1 vssd1 vccd1 vccd1 _09632_/C sky130_fd_sc_hd__nand3_1
XFILLER_56_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09561_ _15650_/Q _09692_/B _09561_/C vssd1 vssd1 vccd1 vccd1 _09561_/X sky130_fd_sc_hd__and3_1
XFILLER_82_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08512_ _08512_/A _08512_/B vssd1 vssd1 vccd1 vccd1 _08512_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09492_ _09507_/C vssd1 vssd1 vccd1 vccd1 _09519_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08443_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08444_/B sky130_fd_sc_hd__xnor2_2
XFILLER_51_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08374_ _08454_/A _08374_/B vssd1 vssd1 vccd1 vccd1 _08374_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09828_ _15701_/Q _10301_/C _09836_/C vssd1 vssd1 vccd1 vccd1 _09828_/Y sky130_fd_sc_hd__nand3_1
XFILLER_47_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09759_ _09770_/C vssd1 vssd1 vccd1 vccd1 _09781_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _16161_/Q _12770_/B _12770_/C vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__and3_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _16012_/Q _11891_/B _11721_/C vssd1 vssd1 vccd1 vccd1 _11731_/A sky130_fd_sc_hd__and3_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14440_ _14441_/B _14441_/C _14387_/X vssd1 vssd1 vccd1 vccd1 _14442_/B sky130_fd_sc_hd__o21ai_1
X_11652_ _11652_/A vssd1 vssd1 vccd1 vccd1 _16001_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ _10649_/A _10603_/B _10603_/C vssd1 vssd1 vccd1 vccd1 _10604_/A sky130_fd_sc_hd__and3_1
X_14371_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14484_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11583_ _11604_/A _11583_/B _11583_/C vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__and3_1
X_16110_ _16118_/CLK _16110_/D vssd1 vssd1 vccd1 vccd1 _16110_/Q sky130_fd_sc_hd__dfxtp_2
X_13322_ _13322_/A vssd1 vssd1 vccd1 vccd1 _13336_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10534_ _15834_/Q _10565_/C _10426_/X vssd1 vssd1 vccd1 vccd1 _10537_/B sky130_fd_sc_hd__a21oi_1
XFILLER_127_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16041_ _16118_/CLK _16041_/D vssd1 vssd1 vccd1 vccd1 _16041_/Q sky130_fd_sc_hd__dfxtp_1
X_10465_ _10465_/A _10465_/B vssd1 vssd1 vccd1 vccd1 _10466_/B sky130_fd_sc_hd__nor2_1
X_13253_ _13249_/Y _13259_/A _13252_/Y _13246_/C vssd1 vssd1 vccd1 vccd1 _13255_/B
+ sky130_fd_sc_hd__o211a_1
X_12204_ _16081_/Q _12204_/B _12204_/C vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__and3_1
XFILLER_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10396_ _15809_/Q _10396_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10396_/Y sky130_fd_sc_hd__nand3_1
X_13184_ _14308_/A vssd1 vssd1 vccd1 vccd1 _13184_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _12304_/A _12135_/B _12135_/C vssd1 vssd1 vccd1 vccd1 _12136_/C sky130_fd_sc_hd__or3_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ _12066_/A _12074_/B vssd1 vssd1 vccd1 vccd1 _12068_/A sky130_fd_sc_hd__or2_1
XFILLER_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11017_ _15913_/Q _11026_/C _10905_/X vssd1 vssd1 vccd1 vccd1 _11017_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15825_ _16595_/CLK _15825_/D vssd1 vssd1 vccd1 vccd1 _15825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15756_ _15812_/CLK _15756_/D vssd1 vssd1 vccd1 vccd1 _15756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ _12968_/A vssd1 vssd1 vccd1 vccd1 _14095_/A sky130_fd_sc_hd__buf_4
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14707_ _14707_/A _14707_/B _14707_/C vssd1 vssd1 vccd1 vccd1 _14708_/A sky130_fd_sc_hd__and3_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11919_ _11940_/A _11919_/B _11919_/C vssd1 vssd1 vccd1 vccd1 _11920_/A sky130_fd_sc_hd__and3_1
X_15687_ _15791_/CLK _15687_/D vssd1 vssd1 vccd1 vccd1 _15687_/Q sky130_fd_sc_hd__dfxtp_1
X_12899_ _12907_/A _12899_/B _12899_/C vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__and3_1
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ _16429_/Q _14640_/C _14411_/X vssd1 vssd1 vccd1 vccd1 _14638_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14569_ _16418_/Q _14569_/B _14576_/C vssd1 vssd1 vccd1 vccd1 _14571_/C sky130_fd_sc_hd__nand3_1
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16308_ _16346_/CLK _16308_/D vssd1 vssd1 vccd1 vccd1 _16308_/Q sky130_fd_sc_hd__dfxtp_1
X_08090_ _08090_/A _08090_/B vssd1 vssd1 vccd1 vccd1 _08276_/B sky130_fd_sc_hd__xor2_1
XFILLER_146_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16239_ _16261_/CLK _16239_/D vssd1 vssd1 vccd1 vccd1 _16239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08992_ _08992_/A _08992_/B vssd1 vssd1 vccd1 vccd1 _08994_/A sky130_fd_sc_hd__or2_1
XFILLER_141_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07943_ _13551_/A _07943_/B vssd1 vssd1 vccd1 vccd1 _07944_/B sky130_fd_sc_hd__xnor2_2
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07874_ _12987_/A _07874_/B vssd1 vssd1 vccd1 vccd1 _07876_/B sky130_fd_sc_hd__xnor2_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09613_ _09438_/X _09611_/B _09530_/X vssd1 vssd1 vccd1 vccd1 _09613_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09544_ _15647_/Q _09585_/B _09550_/C vssd1 vssd1 vccd1 vccd1 _09546_/C sky130_fd_sc_hd__nand3_1
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09475_ _09471_/Y _09474_/X _09431_/X vssd1 vssd1 vccd1 vccd1 _09475_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08426_ _13652_/A vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__clkbuf_2
X_08357_ _08357_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _08357_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08288_ _15624_/Q _08288_/B vssd1 vssd1 vccd1 vccd1 _08288_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10250_ _10250_/A _10250_/B _10250_/C vssd1 vssd1 vccd1 vccd1 _10251_/A sky130_fd_sc_hd__and3_1
XFILLER_106_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ _10486_/A vssd1 vssd1 vccd1 vccd1 _10181_/X sky130_fd_sc_hd__buf_2
XFILLER_121_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _13977_/A _13940_/B _13940_/C vssd1 vssd1 vccd1 vccd1 _13941_/A sky130_fd_sc_hd__and3_1
XFILLER_120_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13871_ _13868_/Y _13877_/A _13870_/Y _13866_/C vssd1 vssd1 vccd1 vccd1 _13873_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15610_ _16551_/CLK _15610_/D vssd1 vssd1 vccd1 vccd1 _15610_/Q sky130_fd_sc_hd__dfxtp_1
X_12822_ _12823_/B _12823_/C _12823_/A vssd1 vssd1 vccd1 vccd1 _12824_/B sky130_fd_sc_hd__a21o_1
X_16590_ _16595_/CLK _16590_/D vssd1 vssd1 vccd1 vccd1 _16590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15541_ _16551_/CLK _15541_/D vssd1 vssd1 vccd1 vccd1 _15541_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12753_ _12868_/A _12753_/B _12753_/C vssd1 vssd1 vccd1 vccd1 _12754_/C sky130_fd_sc_hd__or3_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _12269_/A vssd1 vssd1 vccd1 vccd1 _11928_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15472_ _16570_/CLK _15472_/D vssd1 vssd1 vccd1 vccd1 _15472_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12684_ _16148_/Q _12692_/C _12567_/X vssd1 vssd1 vccd1 vccd1 _12684_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14423_ _14421_/Y _14417_/C _14419_/Y _14420_/X vssd1 vssd1 vccd1 vccd1 _14424_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11635_ _11658_/A _11635_/B _11635_/C vssd1 vssd1 vccd1 vccd1 _11636_/A sky130_fd_sc_hd__and3_1
X_14354_ _14369_/A _14354_/B _14354_/C vssd1 vssd1 vccd1 vccd1 _14355_/A sky130_fd_sc_hd__and3_1
X_11566_ _11619_/A vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ _16236_/Q _13305_/B _13305_/C vssd1 vssd1 vccd1 vccd1 _13313_/A sky130_fd_sc_hd__and3_1
X_10517_ _15830_/Q _10707_/B _10517_/C vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__and3_1
X_14285_ _16375_/Q _14506_/B _14296_/C vssd1 vssd1 vccd1 vccd1 _14291_/A sky130_fd_sc_hd__and3_1
X_11497_ _11495_/Y _11491_/C _11493_/Y _11502_/A vssd1 vssd1 vccd1 vccd1 _11502_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16024_ _16118_/CLK _16024_/D vssd1 vssd1 vccd1 vccd1 _16024_/Q sky130_fd_sc_hd__dfxtp_1
X_13236_ _13233_/Y _13234_/X _13235_/Y _13231_/C vssd1 vssd1 vccd1 vccd1 _13238_/B
+ sky130_fd_sc_hd__o211ai_1
X_10448_ _15818_/Q _10646_/B _10457_/C vssd1 vssd1 vccd1 vccd1 _10448_/Y sky130_fd_sc_hd__nand3_1
XFILLER_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _13190_/A _13167_/B _13167_/C vssd1 vssd1 vccd1 vccd1 _13168_/A sky130_fd_sc_hd__and3_1
X_10379_ _15807_/Q _10483_/B _10379_/C vssd1 vssd1 vccd1 vccd1 _10384_/A sky130_fd_sc_hd__and3_1
X_12118_ _16068_/Q _12173_/B _12118_/C vssd1 vssd1 vccd1 vccd1 _12127_/A sky130_fd_sc_hd__and3_1
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13098_ _13112_/C vssd1 vssd1 vccd1 vccd1 _13120_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12049_ _12049_/A vssd1 vssd1 vccd1 vccd1 _16057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15808_ _15812_/CLK _15808_/D vssd1 vssd1 vccd1 vccd1 _15808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15739_ _15812_/CLK _15739_/D vssd1 vssd1 vccd1 vccd1 _15739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09260_ _09261_/B _09261_/C _09261_/A vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08211_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08212_/B sky130_fd_sc_hd__and2_1
X_09191_ _15578_/Q _09192_/C _10510_/A vssd1 vssd1 vccd1 vccd1 _09193_/A sky130_fd_sc_hd__a21oi_1
X_08142_ _08321_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08143_/B sky130_fd_sc_hd__xor2_1
XFILLER_146_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08073_ _15579_/Q _15561_/Q vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__nand2_1
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08975_ _10430_/A vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__buf_4
XFILLER_103_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07926_ _16598_/Q _16596_/Q vssd1 vssd1 vccd1 vccd1 _07928_/A sky130_fd_sc_hd__or2_1
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07857_ _16514_/Q vssd1 vssd1 vccd1 vccd1 _15069_/A sky130_fd_sc_hd__clkinv_4
XFILLER_84_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07788_ _07806_/A vssd1 vssd1 vccd1 vccd1 _07793_/A sky130_fd_sc_hd__buf_12
X_09527_ _09656_/A _09527_/B vssd1 vssd1 vccd1 vccd1 _09527_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09458_ _15630_/Q _09636_/B _09458_/C vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__and3_1
XFILLER_40_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08409_ _08291_/A _08291_/B _08408_/Y vssd1 vssd1 vccd1 vccd1 _08410_/B sky130_fd_sc_hd__a21oi_1
X_09389_ _15355_/A _09389_/B vssd1 vssd1 vccd1 vccd1 _09390_/B sky130_fd_sc_hd__and2_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ _15969_/Q _11594_/B _11420_/C vssd1 vssd1 vccd1 vccd1 _11420_/Y sky130_fd_sc_hd__nand3_1
XFILLER_61_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11351_ _11351_/A vssd1 vssd1 vccd1 vccd1 _15959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10302_ _10299_/Y _10300_/X _10301_/Y _10297_/C vssd1 vssd1 vccd1 vccd1 _10304_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14070_ _14070_/A vssd1 vssd1 vccd1 vccd1 _16343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ _11850_/A vssd1 vssd1 vccd1 vccd1 _11282_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13021_ _16196_/Q _13028_/C _12850_/X vssd1 vssd1 vccd1 vccd1 _13021_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10233_ _15780_/Q _10267_/C _10176_/X vssd1 vssd1 vccd1 vccd1 _10236_/B sky130_fd_sc_hd__a21oi_1
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10164_ _10414_/A vssd1 vssd1 vccd1 vccd1 _10164_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10095_ _10093_/Y _10089_/C _10091_/Y _10092_/X vssd1 vssd1 vccd1 vccd1 _10096_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14972_ _14972_/A vssd1 vssd1 vccd1 vccd1 _16480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16711_ _16711_/A _07814_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
X_13923_ _16324_/Q _14148_/B _13923_/C vssd1 vssd1 vccd1 vccd1 _13931_/A sky130_fd_sc_hd__and3_1
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13854_ _16314_/Q _13856_/C _13853_/X vssd1 vssd1 vccd1 vccd1 _13854_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_142_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ _13371_/A vssd1 vssd1 vccd1 vccd1 _13034_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16573_ _16595_/CLK _16573_/D vssd1 vssd1 vccd1 vccd1 _16573_/Q sky130_fd_sc_hd__dfxtp_2
X_13785_ _16304_/Q _13793_/C _13729_/X vssd1 vssd1 vccd1 vccd1 _13789_/B sky130_fd_sc_hd__a21o_1
X_10997_ _10995_/A _10995_/B _10996_/X vssd1 vssd1 vccd1 vccd1 _15908_/D sky130_fd_sc_hd__a21oi_1
X_15524_ _16551_/CLK _15524_/D vssd1 vssd1 vccd1 vccd1 _15524_/Q sky130_fd_sc_hd__dfxtp_1
X_12736_ _12736_/A _12736_/B _12736_/C vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__and3_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ _16570_/CLK _15455_/D vssd1 vssd1 vccd1 vccd1 _15455_/Q sky130_fd_sc_hd__dfxtp_2
X_12667_ _12667_/A vssd1 vssd1 vccd1 vccd1 _16144_/D sky130_fd_sc_hd__clkbuf_1
X_14406_ _16393_/Q _14458_/B _14406_/C vssd1 vssd1 vccd1 vccd1 _14406_/X sky130_fd_sc_hd__and3_1
X_11618_ _11616_/A _11616_/B _11617_/X vssd1 vssd1 vccd1 vccd1 _15996_/D sky130_fd_sc_hd__a21oi_1
X_15386_ _15997_/Q _15996_/Q _15995_/Q _15385_/X vssd1 vssd1 vccd1 vccd1 _16570_/D
+ sky130_fd_sc_hd__o31a_1
X_12598_ _13443_/A vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__buf_2
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14337_ _14358_/C vssd1 vssd1 vccd1 vccd1 _14373_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11549_ _11963_/A vssd1 vssd1 vccd1 vccd1 _11666_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14268_ _16373_/Q _14486_/B _14268_/C vssd1 vssd1 vccd1 vccd1 _14276_/B sky130_fd_sc_hd__and3_1
XFILLER_144_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16007_ _16554_/Q _16007_/D vssd1 vssd1 vccd1 vccd1 _16007_/Q sky130_fd_sc_hd__dfxtp_1
X_13219_ _13219_/A _13219_/B _13224_/A vssd1 vssd1 vccd1 vccd1 _16222_/D sky130_fd_sc_hd__nor3_1
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _16364_/Q _14207_/C _13979_/X vssd1 vssd1 vccd1 vccd1 _14199_/Y sky130_fd_sc_hd__a21oi_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08760_ _15485_/Q _08779_/C _08576_/X vssd1 vssd1 vccd1 vccd1 _08762_/B sky130_fd_sc_hd__a21oi_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08691_ _08691_/A _08691_/B vssd1 vssd1 vccd1 vccd1 _08693_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09312_ _09749_/A _10526_/A _09296_/B _08554_/A vssd1 vssd1 vccd1 vccd1 _09313_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09243_ _09243_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _15585_/D sky130_fd_sc_hd__nor2_1
X_09174_ _15575_/Q _15332_/B _09178_/C vssd1 vssd1 vccd1 vccd1 _09180_/A sky130_fd_sc_hd__and3_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08125_ _07892_/A _07892_/B _08124_/Y vssd1 vssd1 vccd1 vccd1 _08137_/A sky130_fd_sc_hd__o21ai_4
XFILLER_147_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08056_ _15687_/Q _15669_/Q vssd1 vssd1 vccd1 vccd1 _08058_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08958_ _09037_/A _08963_/C vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__and2_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07909_ _16610_/Q _16608_/Q vssd1 vssd1 vccd1 vccd1 _07910_/B sky130_fd_sc_hd__or2_1
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08889_ _15525_/Q vssd1 vssd1 vccd1 vccd1 _08896_/C sky130_fd_sc_hd__inv_2
XFILLER_57_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10920_ _15899_/Q _10928_/C _10919_/X vssd1 vssd1 vccd1 vccd1 _10920_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16680__85 vssd1 vssd1 vccd1 vccd1 _16680__85/HI _16756_/A sky130_fd_sc_hd__conb_1
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ _15890_/Q _11076_/B _10852_/C vssd1 vssd1 vccd1 vccd1 _10851_/X sky130_fd_sc_hd__and3_1
XFILLER_72_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _14411_/A vssd1 vssd1 vccd1 vccd1 _13570_/X sky130_fd_sc_hd__clkbuf_2
X_10782_ _15880_/Q _10782_/B _10782_/C vssd1 vssd1 vccd1 vccd1 _10782_/X sky130_fd_sc_hd__and3_1
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12749_/A _12526_/C vssd1 vssd1 vccd1 vccd1 _12521_/X sky130_fd_sc_hd__or2_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _16527_/Q _15248_/C _10782_/B vssd1 vssd1 vccd1 vccd1 _15240_/Y sky130_fd_sc_hd__a21oi_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _12450_/Y _12446_/C _12448_/Y _12449_/X vssd1 vssd1 vccd1 vccd1 _12453_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11403_ _11520_/A _11403_/B _11407_/A vssd1 vssd1 vccd1 vccd1 _15966_/D sky130_fd_sc_hd__nor3_1
X_15171_ _15171_/A vssd1 vssd1 vccd1 vccd1 _16513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12383_ _12398_/A _12383_/B _12383_/C vssd1 vssd1 vccd1 vccd1 _12384_/A sky130_fd_sc_hd__and3_1
XFILLER_125_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ _14123_/B _14123_/C _14123_/A vssd1 vssd1 vccd1 vccd1 _14124_/B sky130_fd_sc_hd__a21o_1
X_11334_ _11334_/A vssd1 vssd1 vccd1 vccd1 _11371_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14053_ _14276_/A _14053_/B _14053_/C vssd1 vssd1 vccd1 vccd1 _14054_/C sky130_fd_sc_hd__or3_1
X_11265_ _11265_/A vssd1 vssd1 vccd1 vccd1 _15946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13004_ _13019_/A _13004_/B _13004_/C vssd1 vssd1 vccd1 vccd1 _13005_/A sky130_fd_sc_hd__and3_1
X_10216_ _10216_/A _10216_/B vssd1 vssd1 vccd1 vccd1 _10217_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11196_ _15938_/Q _11359_/B _11197_/C vssd1 vssd1 vccd1 vccd1 _11196_/X sky130_fd_sc_hd__and3_1
XFILLER_97_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _15766_/Q _10158_/C _10009_/B vssd1 vssd1 vccd1 vccd1 _10147_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14955_ _14956_/B _14956_/C _14954_/X vssd1 vssd1 vccd1 vccd1 _14957_/B sky130_fd_sc_hd__o21ai_1
X_10078_ _15754_/Q _10086_/C _10729_/B vssd1 vssd1 vccd1 vccd1 _10081_/B sky130_fd_sc_hd__a21o_1
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13906_ _16322_/Q _13906_/B _13908_/C vssd1 vssd1 vccd1 vccd1 _13906_/X sky130_fd_sc_hd__and3_1
X_14886_ _16468_/Q _14887_/C _14828_/X vssd1 vssd1 vccd1 vccd1 _14888_/A sky130_fd_sc_hd__a21oi_1
XFILLER_62_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13837_ _13869_/C vssd1 vssd1 vccd1 vccd1 _13875_/C sky130_fd_sc_hd__clkbuf_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16556_ _16570_/CLK _16556_/D vssd1 vssd1 vccd1 vccd1 _16556_/Q sky130_fd_sc_hd__dfxtp_1
X_13768_ _13768_/A _13768_/B vssd1 vssd1 vccd1 vccd1 _13774_/C sky130_fd_sc_hd__nor2_1
XFILLER_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12719_ _12717_/Y _12718_/X _12714_/C _12715_/C vssd1 vssd1 vccd1 vccd1 _12721_/B
+ sky130_fd_sc_hd__o211ai_1
X_15507_ _16551_/CLK _15507_/D vssd1 vssd1 vccd1 vccd1 _15507_/Q sky130_fd_sc_hd__dfxtp_1
X_16487_ _16607_/CLK _16487_/D vssd1 vssd1 vccd1 vccd1 _16487_/Q sky130_fd_sc_hd__dfxtp_1
X_13699_ _16292_/Q _13709_/C _13698_/X vssd1 vssd1 vccd1 vccd1 _13699_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15438_ _16339_/Q _16341_/Q _16340_/Q _15434_/X vssd1 vssd1 vccd1 vccd1 _16613_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _15893_/Q _15892_/Q _15891_/Q _15363_/X vssd1 vssd1 vccd1 vccd1 _16557_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_116_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09930_ _09924_/Y _09925_/X _09927_/B vssd1 vssd1 vccd1 vccd1 _09931_/B sky130_fd_sc_hd__o21a_1
XFILLER_131_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09861_ _09864_/C vssd1 vssd1 vccd1 vccd1 _09873_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08812_ _15496_/Q _08822_/C _08604_/X vssd1 vssd1 vccd1 vccd1 _08812_/Y sky130_fd_sc_hd__a21oi_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09792_ _09792_/A vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__clkbuf_2
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08831_/A _08752_/C vssd1 vssd1 vccd1 vccd1 _08745_/A sky130_fd_sc_hd__and2_1
XFILLER_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08674_ _10285_/C vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__buf_2
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09226_ _15586_/Q _15341_/B _09231_/C vssd1 vssd1 vccd1 vccd1 _09233_/A sky130_fd_sc_hd__and3_1
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09157_ _09151_/B _09154_/B _09117_/X vssd1 vssd1 vccd1 vccd1 _09165_/C sky130_fd_sc_hd__o21a_1
XFILLER_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08108_ _08108_/A _16703_/A _15282_/C vssd1 vssd1 vccd1 vccd1 _08109_/C sky130_fd_sc_hd__nor3_1
X_09088_ _09006_/X _09086_/A _08927_/X vssd1 vssd1 vccd1 vccd1 _09088_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08039_ _08039_/A _08039_/B vssd1 vssd1 vccd1 vccd1 _08051_/A sky130_fd_sc_hd__and2_4
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11050_ _11048_/A _11048_/B _11049_/X vssd1 vssd1 vccd1 vccd1 _15916_/D sky130_fd_sc_hd__a21oi_1
XFILLER_131_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10001_ _10055_/A _10001_/B _10004_/B vssd1 vssd1 vccd1 vccd1 _15735_/D sky130_fd_sc_hd__nor3_1
XFILLER_77_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14740_ _14740_/A vssd1 vssd1 vccd1 vccd1 _16444_/D sky130_fd_sc_hd__clkbuf_1
X_11952_ _11952_/A _11952_/B vssd1 vssd1 vccd1 vccd1 _11954_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _10925_/A _10903_/B _10903_/C vssd1 vssd1 vccd1 vccd1 _10904_/A sky130_fd_sc_hd__and3_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14671_ _14839_/A _14671_/B _14671_/C vssd1 vssd1 vccd1 vccd1 _14672_/C sky130_fd_sc_hd__or3_1
X_11883_ _16035_/Q _11891_/C _11770_/X vssd1 vssd1 vccd1 vccd1 _11883_/Y sky130_fd_sc_hd__a21oi_1
X_16410_ input11/X _16410_/D vssd1 vssd1 vccd1 vccd1 _16410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13622_ _16282_/Q _13625_/C _13570_/X vssd1 vssd1 vccd1 vccd1 _13622_/Y sky130_fd_sc_hd__a21oi_1
X_10834_ _10954_/A _10834_/B _10838_/A vssd1 vssd1 vccd1 vccd1 _15886_/D sky130_fd_sc_hd__nor3_1
Xrepeater13 _16553_/Q vssd1 vssd1 vccd1 vccd1 _15365_/A sky130_fd_sc_hd__buf_12
Xrepeater24 input11/X vssd1 vssd1 vccd1 vccd1 _15812_/CLK sky130_fd_sc_hd__buf_12
X_16341_ _16346_/CLK _16341_/D vssd1 vssd1 vccd1 vccd1 _16341_/Q sky130_fd_sc_hd__dfxtp_1
X_13553_ _13573_/C vssd1 vssd1 vccd1 vccd1 _13586_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10765_ _08663_/X _10762_/B _10764_/Y vssd1 vssd1 vccd1 vccd1 _15875_/D sky130_fd_sc_hd__o21a_1
X_12504_ _12502_/Y _12498_/C _12500_/Y _12501_/X vssd1 vssd1 vccd1 vccd1 _12505_/C
+ sky130_fd_sc_hd__a211o_1
X_16272_ _16533_/Q _16272_/D vssd1 vssd1 vccd1 vccd1 _16272_/Q sky130_fd_sc_hd__dfxtp_1
X_13484_ _13482_/A _13482_/B _13483_/X vssd1 vssd1 vccd1 vccd1 _16260_/D sky130_fd_sc_hd__a21oi_1
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10696_ _10696_/A vssd1 vssd1 vccd1 vccd1 _15862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15223_ _15274_/A _15223_/B _15223_/C vssd1 vssd1 vccd1 vccd1 _15224_/C sky130_fd_sc_hd__or3_1
XFILLER_32_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ _16113_/Q _12487_/B _12435_/C vssd1 vssd1 vccd1 vccd1 _12435_/X sky130_fd_sc_hd__and3_1
XFILLER_32_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15154_ _16512_/Q _15161_/C _08747_/A vssd1 vssd1 vccd1 vccd1 _15154_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12366_ _12387_/C vssd1 vssd1 vccd1 vccd1 _12402_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ _14158_/A _14110_/C vssd1 vssd1 vccd1 vccd1 _14105_/X sky130_fd_sc_hd__or2_1
X_11317_ _11314_/Y _11315_/X _11316_/Y _11312_/C vssd1 vssd1 vccd1 vccd1 _11319_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15085_ _15079_/C _15080_/C _15082_/Y _15083_/X vssd1 vssd1 vccd1 vccd1 _15086_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12297_ _12297_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12299_/A sky130_fd_sc_hd__or2_1
XFILLER_4_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14036_ _14036_/A vssd1 vssd1 vccd1 vccd1 _16338_/D sky130_fd_sc_hd__clkbuf_1
X_11248_ _11242_/C _11243_/C _11245_/Y _11246_/X vssd1 vssd1 vccd1 vccd1 _11249_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_121_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11179_ _15935_/Q _11402_/B _11190_/C vssd1 vssd1 vccd1 vccd1 _11185_/A sky130_fd_sc_hd__and3_1
XFILLER_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15987_ _16005_/CLK _15987_/D vssd1 vssd1 vccd1 vccd1 _15987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14938_ _15207_/A vssd1 vssd1 vccd1 vccd1 _15053_/A sky130_fd_sc_hd__buf_2
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14869_ _14867_/Y _14863_/C _14865_/Y _14866_/X vssd1 vssd1 vccd1 vccd1 _14870_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16608_ input11/X _16608_/D vssd1 vssd1 vccd1 vccd1 _16608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08390_ _08458_/A _08458_/B vssd1 vssd1 vccd1 vccd1 _08393_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16539_ _16595_/CLK _16539_/D vssd1 vssd1 vccd1 vccd1 _16708_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09011_ _15539_/Q _09028_/C _08843_/X vssd1 vssd1 vccd1 vccd1 _09013_/B sky130_fd_sc_hd__a21oi_1
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09913_ _15720_/Q _09914_/C _08604_/A vssd1 vssd1 vccd1 vccd1 _09913_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _11150_/A vssd1 vssd1 vccd1 vccd1 _10313_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _15694_/Q _09919_/B _09781_/C vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__and3_1
XFILLER_74_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08726_ _15478_/Q _08732_/C _08604_/X vssd1 vssd1 vccd1 vccd1 _08726_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ input7/X vssd1 vssd1 vccd1 vccd1 _14895_/A sky130_fd_sc_hd__buf_2
XFILLER_82_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16650__55 vssd1 vssd1 vccd1 vccd1 _16650__55/HI _16726_/A sky130_fd_sc_hd__conb_1
XFILLER_42_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08588_ _10183_/A vssd1 vssd1 vccd1 vccd1 _08589_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ _10550_/A vssd1 vssd1 vccd1 vccd1 _15834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09209_ _09087_/X _09206_/A _09208_/Y vssd1 vssd1 vccd1 vccd1 _15578_/D sky130_fd_sc_hd__o21a_1
XFILLER_10_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10481_ _10509_/C vssd1 vssd1 vccd1 vccd1 _10517_/C sky130_fd_sc_hd__clkbuf_2
X_12220_ _12217_/Y _12218_/X _12219_/Y _12215_/C vssd1 vssd1 vccd1 vccd1 _12222_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12151_ _16073_/Q _12160_/C _12036_/X vssd1 vssd1 vccd1 vccd1 _12151_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11102_ _11384_/A vssd1 vssd1 vccd1 vccd1 _11332_/A sky130_fd_sc_hd__buf_2
X_12082_ _16063_/Q _12125_/C _12081_/X vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11033_ _15914_/Q _11205_/B _11039_/C vssd1 vssd1 vccd1 vccd1 _11033_/Y sky130_fd_sc_hd__nand3_1
X_15910_ _16553_/Q _15910_/D vssd1 vssd1 vccd1 vccd1 _15910_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15841_ _16595_/CLK _15841_/D vssd1 vssd1 vccd1 vccd1 _15841_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15772_ _15791_/CLK _15772_/D vssd1 vssd1 vccd1 vccd1 _15772_/Q sky130_fd_sc_hd__dfxtp_1
X_12984_ _13151_/A _12984_/B _12984_/C vssd1 vssd1 vccd1 vccd1 _12985_/C sky130_fd_sc_hd__or3_1
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14723_ _14724_/B _14724_/C _14669_/X vssd1 vssd1 vccd1 vccd1 _14725_/B sky130_fd_sc_hd__o21ai_1
X_11935_ _16043_/Q _11944_/C _11770_/X vssd1 vssd1 vccd1 vccd1 _11935_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14654_ _16431_/Q _14662_/C _14537_/X vssd1 vssd1 vccd1 vccd1 _14654_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11866_ _11888_/A _11866_/B _11866_/C vssd1 vssd1 vccd1 vccd1 _11867_/A sky130_fd_sc_hd__and3_1
X_13605_ _13625_/C vssd1 vssd1 vccd1 vccd1 _13639_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10817_ _11049_/A _10823_/C vssd1 vssd1 vccd1 vccd1 _10817_/X sky130_fd_sc_hd__or2_1
X_14585_ _14583_/Y _14579_/C _14581_/Y _14582_/X vssd1 vssd1 vccd1 vccd1 _14586_/C
+ sky130_fd_sc_hd__a211o_1
X_11797_ _11797_/A vssd1 vssd1 vccd1 vccd1 _16021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13536_ _13643_/A _13536_/B _13540_/B vssd1 vssd1 vccd1 vccd1 _16267_/D sky130_fd_sc_hd__nor3_1
X_16324_ _16346_/CLK _16324_/D vssd1 vssd1 vccd1 vccd1 _16324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10748_ _15874_/Q _10755_/C _09604_/A vssd1 vssd1 vccd1 vccd1 _10748_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16255_ _16261_/CLK _16255_/D vssd1 vssd1 vccd1 vccd1 _16255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13467_ _16258_/Q _13467_/B _13473_/C vssd1 vssd1 vccd1 vccd1 _13467_/Y sky130_fd_sc_hd__nand3_1
X_10679_ _15862_/Q _10679_/B _10685_/C vssd1 vssd1 vccd1 vccd1 _10681_/C sky130_fd_sc_hd__nand3_1
X_15206_ _15206_/A vssd1 vssd1 vccd1 vccd1 _16519_/D sky130_fd_sc_hd__clkbuf_1
X_12418_ _12586_/A _12418_/B _12418_/C vssd1 vssd1 vccd1 vccd1 _12419_/C sky130_fd_sc_hd__or3_1
X_16186_ _16237_/CLK _16186_/D vssd1 vssd1 vccd1 vccd1 _16186_/Q sky130_fd_sc_hd__dfxtp_1
X_13398_ _16250_/Q _13401_/C _13289_/X vssd1 vssd1 vccd1 vccd1 _13398_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ _15131_/C _15132_/C _15134_/Y _15135_/X vssd1 vssd1 vccd1 vccd1 _15138_/C
+ sky130_fd_sc_hd__a211o_1
X_12349_ _12347_/Y _12343_/C _12345_/Y _12354_/A vssd1 vssd1 vccd1 vccd1 _12354_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15068_ _15207_/A vssd1 vssd1 vccd1 vccd1 _15180_/A sky130_fd_sc_hd__buf_2
XFILLER_142_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14019_ _14012_/C _14013_/C _14016_/Y _14017_/X vssd1 vssd1 vccd1 vccd1 _14020_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07890_ _08132_/A _08132_/B vssd1 vssd1 vccd1 vccd1 _08124_/B sky130_fd_sc_hd__xor2_4
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _09557_/A _09556_/Y _09557_/B vssd1 vssd1 vccd1 vccd1 _09560_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08511_ _08537_/A _08537_/B vssd1 vssd1 vccd1 vccd1 _08535_/A sky130_fd_sc_hd__xnor2_4
XFILLER_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09491_ _09496_/C vssd1 vssd1 vccd1 vccd1 _09507_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08442_ _08351_/A _08351_/B _08353_/B _08353_/A vssd1 vssd1 vccd1 vccd1 _08443_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_91_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08373_ _08454_/B _08373_/B vssd1 vssd1 vccd1 vccd1 _08374_/B sky130_fd_sc_hd__and2b_1
XFILLER_32_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09827_ _10447_/A vssd1 vssd1 vccd1 vccd1 _10301_/C sky130_fd_sc_hd__buf_4
XFILLER_74_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09758_ _09761_/C vssd1 vssd1 vccd1 vccd1 _09770_/C sky130_fd_sc_hd__clkbuf_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ _08706_/X _08704_/A _08708_/X vssd1 vssd1 vccd1 vccd1 _08710_/B sky130_fd_sc_hd__o21ai_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _09688_/X _09687_/Y _09644_/X vssd1 vssd1 vccd1 vccd1 _09689_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _16012_/Q _11729_/C _11719_/X vssd1 vssd1 vccd1 vccd1 _11720_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11651_ _11658_/A _11651_/B _11651_/C vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__and3_1
XFILLER_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10602_ _10600_/Y _10596_/C _10598_/Y _10599_/X vssd1 vssd1 vccd1 vccd1 _10603_/C
+ sky130_fd_sc_hd__a211o_1
X_14370_ _14370_/A vssd1 vssd1 vccd1 vccd1 _16386_/D sky130_fd_sc_hd__clkbuf_1
X_11582_ _11582_/A _11582_/B _11582_/C vssd1 vssd1 vccd1 vccd1 _11583_/C sky130_fd_sc_hd__nand3_1
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13321_ _13321_/A vssd1 vssd1 vccd1 vccd1 _16237_/D sky130_fd_sc_hd__clkbuf_1
X_10533_ _10559_/C vssd1 vssd1 vccd1 vccd1 _10565_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16040_ _16118_/CLK _16040_/D vssd1 vssd1 vccd1 vccd1 _16040_/Q sky130_fd_sc_hd__dfxtp_1
X_13252_ _16227_/Q _13474_/B _13257_/C vssd1 vssd1 vccd1 vccd1 _13252_/Y sky130_fd_sc_hd__nand3_1
X_10464_ _10464_/A _10464_/B vssd1 vssd1 vccd1 vccd1 _10466_/A sky130_fd_sc_hd__or2_1
XFILLER_89_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12203_ _16081_/Q _12212_/C _12036_/X vssd1 vssd1 vccd1 vccd1 _12203_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13183_ _13183_/A vssd1 vssd1 vccd1 vccd1 _14308_/A sky130_fd_sc_hd__buf_4
X_10395_ _15810_/Q _10446_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__and3_1
XFILLER_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12134_ _12135_/B _12135_/C _12133_/X vssd1 vssd1 vccd1 vccd1 _12136_/B sky130_fd_sc_hd__o21ai_1
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12065_ _16061_/Q _12232_/B _12065_/C vssd1 vssd1 vccd1 vccd1 _12074_/B sky130_fd_sc_hd__and3_1
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11016_ _11016_/A vssd1 vssd1 vccd1 vccd1 _15911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15824_ _16595_/CLK _15824_/D vssd1 vssd1 vccd1 vccd1 _15824_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15755_ _15791_/CLK _15755_/D vssd1 vssd1 vccd1 vccd1 _15755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12967_ _16188_/Q _13022_/B _12967_/C vssd1 vssd1 vccd1 vccd1 _12977_/A sky130_fd_sc_hd__and3_1
X_14706_ _14704_/Y _14700_/C _14702_/Y _14703_/X vssd1 vssd1 vccd1 vccd1 _14707_/C
+ sky130_fd_sc_hd__a211o_1
X_11918_ _11918_/A _11918_/B _11918_/C vssd1 vssd1 vccd1 vccd1 _11919_/C sky130_fd_sc_hd__nand3_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15686_ _15791_/CLK _15686_/D vssd1 vssd1 vccd1 vccd1 _15686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12898_ _12896_/Y _12892_/C _12894_/Y _12895_/X vssd1 vssd1 vccd1 vccd1 _12899_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11849_ _11903_/A vssd1 vssd1 vccd1 vccd1 _11888_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14637_ _14637_/A vssd1 vssd1 vccd1 vccd1 _16427_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _16418_/Q _14576_/C _14567_/X vssd1 vssd1 vccd1 vccd1 _14571_/B sky130_fd_sc_hd__a21o_1
XFILLER_119_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16307_ _16346_/CLK _16307_/D vssd1 vssd1 vccd1 vccd1 _16307_/Q sky130_fd_sc_hd__dfxtp_1
X_13519_ _16267_/Q _13531_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13519_/Y sky130_fd_sc_hd__a21oi_1
X_14499_ _16531_/Q _16530_/Q _16529_/Q _10719_/X vssd1 vssd1 vccd1 vccd1 _16406_/D
+ sky130_fd_sc_hd__o31a_1
X_16238_ _16261_/CLK _16238_/D vssd1 vssd1 vccd1 vccd1 _16238_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_134_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16169_ _16237_/CLK _16169_/D vssd1 vssd1 vccd1 vccd1 _16169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08991_ _15533_/Q _08991_/B _08991_/C vssd1 vssd1 vccd1 vccd1 _08992_/B sky130_fd_sc_hd__and3_1
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07942_ _16607_/Q _08167_/B vssd1 vssd1 vccd1 vccd1 _07943_/B sky130_fd_sc_hd__xnor2_1
XFILLER_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07873_ _14960_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07874_/B sky130_fd_sc_hd__xnor2_4
X_09612_ _09524_/X _09610_/B _09611_/Y vssd1 vssd1 vccd1 vccd1 _15657_/D sky130_fd_sc_hd__o21a_1
XFILLER_83_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09543_ _15647_/Q _09550_/C _09362_/X vssd1 vssd1 vccd1 vccd1 _09546_/B sky130_fd_sc_hd__a21o_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09474_ _09472_/X _09474_/B vssd1 vssd1 vccd1 vccd1 _09474_/X sky130_fd_sc_hd__and2b_1
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16620__25 vssd1 vssd1 vccd1 vccd1 _16620__25/HI _16686_/A sky130_fd_sc_hd__conb_1
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08425_ _08526_/A vssd1 vssd1 vccd1 vccd1 _13652_/A sky130_fd_sc_hd__buf_6
XFILLER_52_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08356_ _08357_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _08356_/X sky130_fd_sc_hd__and2_1
XFILLER_149_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08287_ _08287_/A _08287_/B vssd1 vssd1 vccd1 vccd1 _08408_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10180_ _10340_/A vssd1 vssd1 vccd1 vccd1 _10250_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13870_ _16315_/Q _14039_/B _13875_/C vssd1 vssd1 vccd1 vccd1 _13870_/Y sky130_fd_sc_hd__nand3_1
XFILLER_75_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12821_ _16168_/Q _12881_/B _12828_/C vssd1 vssd1 vccd1 vccd1 _12823_/C sky130_fd_sc_hd__nand3_1
XFILLER_43_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15540_ _16551_/CLK _15540_/D vssd1 vssd1 vccd1 vccd1 _15540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _12753_/B _12753_/C _12699_/X vssd1 vssd1 vccd1 vccd1 _12754_/B sky130_fd_sc_hd__o21ai_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11703_ _16010_/Q _11706_/C _11591_/X vssd1 vssd1 vccd1 vccd1 _11703_/Y sky130_fd_sc_hd__a21oi_1
X_15471_ _16551_/CLK _15471_/D vssd1 vssd1 vccd1 vccd1 _15471_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12683_/A vssd1 vssd1 vccd1 vccd1 _12796_/A sky130_fd_sc_hd__buf_2
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14419_/Y _14420_/X _14421_/Y _14417_/C vssd1 vssd1 vccd1 vccd1 _14424_/B
+ sky130_fd_sc_hd__o211ai_1
X_11634_ _11634_/A _11634_/B _11634_/C vssd1 vssd1 vccd1 vccd1 _11635_/C sky130_fd_sc_hd__nand3_1
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _14347_/C _14348_/C _14350_/Y _14351_/X vssd1 vssd1 vccd1 vccd1 _14354_/C
+ sky130_fd_sc_hd__a211o_1
X_11565_ _11563_/A _11563_/B _11564_/X vssd1 vssd1 vccd1 vccd1 _15988_/D sky130_fd_sc_hd__a21oi_1
X_13304_ _16236_/Q _13311_/C _13133_/X vssd1 vssd1 vccd1 vccd1 _13304_/Y sky130_fd_sc_hd__a21oi_1
X_10516_ _11150_/A vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14284_ _14848_/A vssd1 vssd1 vccd1 vccd1 _14506_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11496_ _11493_/Y _11502_/A _11495_/Y _11491_/C vssd1 vssd1 vccd1 vccd1 _11498_/B
+ sky130_fd_sc_hd__o211a_1
X_16023_ _16118_/CLK _16023_/D vssd1 vssd1 vccd1 vccd1 _16023_/Q sky130_fd_sc_hd__dfxtp_1
X_13235_ _16225_/Q _13292_/B _13235_/C vssd1 vssd1 vccd1 vccd1 _13235_/Y sky130_fd_sc_hd__nand3_1
XFILLER_6_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10447_ _10447_/A vssd1 vssd1 vccd1 vccd1 _10646_/B sky130_fd_sc_hd__clkbuf_2
X_13166_ _13166_/A _13166_/B _13166_/C vssd1 vssd1 vccd1 vccd1 _13167_/C sky130_fd_sc_hd__nand3_1
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10378_ _15807_/Q _10408_/C _10176_/X vssd1 vssd1 vccd1 vccd1 _10380_/B sky130_fd_sc_hd__a21oi_1
XFILLER_112_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12117_ _16068_/Q _12125_/C _12000_/X vssd1 vssd1 vccd1 vccd1 _12117_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13097_ _13097_/A vssd1 vssd1 vccd1 vccd1 _13112_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12048_ _12056_/A _12048_/B _12048_/C vssd1 vssd1 vccd1 vccd1 _12049_/A sky130_fd_sc_hd__and3_1
XFILLER_111_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15807_ _16595_/CLK _15807_/D vssd1 vssd1 vccd1 vccd1 _15807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13999_ _13999_/A vssd1 vssd1 vccd1 vccd1 _16333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15738_ _16551_/CLK _15738_/D vssd1 vssd1 vccd1 vccd1 _15738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15669_ _15791_/CLK _15669_/D vssd1 vssd1 vccd1 vccd1 _15669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08210_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09190_ _10922_/B vssd1 vssd1 vccd1 vccd1 _10510_/A sky130_fd_sc_hd__clkbuf_4
X_08141_ _09255_/C _07896_/B _08140_/X vssd1 vssd1 vccd1 vccd1 _08321_/B sky130_fd_sc_hd__o21a_1
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _15597_/Q vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__clkinv_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08974_ _09054_/A _08974_/B _08980_/A vssd1 vssd1 vccd1 vccd1 _15526_/D sky130_fd_sc_hd__nor3_1
XFILLER_102_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07925_ _16600_/Q vssd1 vssd1 vccd1 vccd1 _13269_/A sky130_fd_sc_hd__clkinv_2
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07856_ _15498_/Q vssd1 vssd1 vccd1 vccd1 _08110_/A sky130_fd_sc_hd__inv_2
XFILLER_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07787_ _07787_/A vssd1 vssd1 vccd1 vccd1 _07787_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09526_ _09655_/A _09526_/B vssd1 vssd1 vccd1 vccd1 _09527_/B sky130_fd_sc_hd__and2_1
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09457_ _10492_/A vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08408_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08408_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09388_ _09381_/Y _09382_/X _09385_/B vssd1 vssd1 vccd1 vccd1 _09389_/B sky130_fd_sc_hd__o21a_1
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08339_ _08339_/A _08440_/A vssd1 vssd1 vccd1 vccd1 _08435_/A sky130_fd_sc_hd__xor2_4
XFILLER_138_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11350_ _11371_/A _11350_/B _11350_/C vssd1 vssd1 vccd1 vccd1 _11351_/A sky130_fd_sc_hd__and3_1
XFILLER_137_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10301_ _15791_/Q _10307_/B _10301_/C vssd1 vssd1 vccd1 vccd1 _10301_/Y sky130_fd_sc_hd__nand3_1
X_11281_ _11334_/A vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13020_ _13020_/A vssd1 vssd1 vccd1 vccd1 _16194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10232_ _10261_/C vssd1 vssd1 vccd1 vccd1 _10267_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_121_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10163_ _10161_/A _10161_/B _10162_/X vssd1 vssd1 vccd1 vccd1 _15765_/D sky130_fd_sc_hd__a21oi_1
XFILLER_120_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10094_ _10091_/Y _10092_/X _10093_/Y _10089_/C vssd1 vssd1 vccd1 vccd1 _10096_/B
+ sky130_fd_sc_hd__o211ai_1
X_14971_ _14992_/A _14971_/B _14971_/C vssd1 vssd1 vccd1 vccd1 _14972_/A sky130_fd_sc_hd__and3_1
XFILLER_120_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16710_ _16710_/A _07811_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13922_ _15048_/A vssd1 vssd1 vccd1 vccd1 _14148_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13853_ _14411_/A vssd1 vssd1 vccd1 vccd1 _13853_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ _12802_/A _12802_/B _12803_/X vssd1 vssd1 vccd1 vccd1 _16164_/D sky130_fd_sc_hd__a21oi_1
X_16572_ _16595_/CLK _16572_/D vssd1 vssd1 vccd1 vccd1 _16572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13784_ _13784_/A _13784_/B _13789_/A vssd1 vssd1 vccd1 vccd1 _16302_/D sky130_fd_sc_hd__nor3_1
X_10996_ _11049_/A _11001_/C vssd1 vssd1 vccd1 vccd1 _10996_/X sky130_fd_sc_hd__or2_1
X_15523_ _16551_/CLK _15523_/D vssd1 vssd1 vccd1 vccd1 _15523_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12733_/Y _12729_/C _12731_/Y _12732_/X vssd1 vssd1 vccd1 vccd1 _12736_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12681_/A _12666_/B _12666_/C vssd1 vssd1 vccd1 vccd1 _12667_/A sky130_fd_sc_hd__and3_1
X_15454_ _16570_/CLK _15454_/D vssd1 vssd1 vccd1 vccd1 _15454_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ _11617_/A _11621_/C vssd1 vssd1 vccd1 vccd1 _11617_/X sky130_fd_sc_hd__or2_1
X_14405_ _16393_/Q _14414_/C _14294_/X vssd1 vssd1 vccd1 vccd1 _14405_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12597_ _12653_/A _12597_/B _12602_/A vssd1 vssd1 vccd1 vccd1 _16134_/D sky130_fd_sc_hd__nor3_1
X_15385_ _15409_/A vssd1 vssd1 vccd1 vccd1 _15385_/X sky130_fd_sc_hd__buf_2
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11548_ _11548_/A vssd1 vssd1 vccd1 vccd1 _15986_/D sky130_fd_sc_hd__clkbuf_1
X_14336_ _14351_/C vssd1 vssd1 vccd1 vccd1 _14358_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14267_ _14830_/A vssd1 vssd1 vccd1 vccd1 _14486_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_11479_ _15978_/Q _11644_/B _11480_/C vssd1 vssd1 vccd1 vccd1 _11479_/X sky130_fd_sc_hd__and3_1
X_13218_ _16223_/Q _13383_/B _13228_/C vssd1 vssd1 vccd1 vccd1 _13224_/A sky130_fd_sc_hd__and3_1
XFILLER_143_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16006_ _16554_/Q _16006_/D vssd1 vssd1 vccd1 vccd1 _16006_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14198_ _14198_/A vssd1 vssd1 vccd1 vccd1 _16362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13317_/A vssd1 vssd1 vccd1 vccd1 _13190_/A sky130_fd_sc_hd__clkbuf_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08690_ _08690_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _08693_/A sky130_fd_sc_hd__or2_1
XFILLER_53_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09311_ _11850_/A vssd1 vssd1 vccd1 vccd1 _10526_/A sky130_fd_sc_hd__buf_2
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09242_ _09744_/A _09244_/C _08667_/A vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09173_ _15575_/Q _09192_/C _09051_/X vssd1 vssd1 vccd1 vccd1 _09175_/B sky130_fd_sc_hd__a21oi_1
XFILLER_119_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08124_ _16568_/Q _08124_/B vssd1 vssd1 vccd1 vccd1 _08124_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08055_ _15705_/Q vssd1 vssd1 vccd1 vccd1 _09761_/C sky130_fd_sc_hd__clkinv_2
XFILLER_135_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08957_ _08872_/X _08949_/B _08952_/B _08956_/Y vssd1 vssd1 vccd1 vccd1 _15521_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07908_ _16610_/Q _16608_/Q vssd1 vssd1 vccd1 vccd1 _07910_/A sky130_fd_sc_hd__nand2_1
X_08888_ _15497_/Q _15496_/Q _15495_/Q _08887_/X vssd1 vssd1 vccd1 vccd1 _15507_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07839_ _07842_/A vssd1 vssd1 vccd1 vccd1 _07839_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10850_ _14979_/A vssd1 vssd1 vccd1 vccd1 _11076_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09509_ _09501_/C _09502_/C _09506_/Y _09513_/A vssd1 vssd1 vccd1 vccd1 _09513_/B
+ sky130_fd_sc_hd__a211oi_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _15880_/Q _10791_/C _15034_/A vssd1 vssd1 vccd1 vccd1 _10781_/Y sky130_fd_sc_hd__a21oi_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12520_/A _12520_/B vssd1 vssd1 vccd1 vccd1 _12526_/C sky130_fd_sc_hd__nor2_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12448_/Y _12449_/X _12450_/Y _12446_/C vssd1 vssd1 vccd1 vccd1 _12453_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11402_ _15967_/Q _11402_/B _11412_/C vssd1 vssd1 vccd1 vccd1 _11407_/A sky130_fd_sc_hd__and3_1
X_15170_ _15205_/A _15170_/B _15170_/C vssd1 vssd1 vccd1 vccd1 _15171_/A sky130_fd_sc_hd__and3_1
X_12382_ _12376_/C _12377_/C _12379_/Y _12380_/X vssd1 vssd1 vccd1 vccd1 _12383_/C
+ sky130_fd_sc_hd__a211o_1
X_14121_ _16352_/Q _14289_/B _14127_/C vssd1 vssd1 vccd1 vccd1 _14123_/C sky130_fd_sc_hd__nand3_1
X_11333_ _11331_/A _11331_/B _11332_/X vssd1 vssd1 vccd1 vccd1 _15956_/D sky130_fd_sc_hd__a21oi_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14052_ _14331_/A vssd1 vssd1 vccd1 vccd1 _14276_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11264_ _11264_/A _11264_/B _11264_/C vssd1 vssd1 vccd1 vccd1 _11265_/A sky130_fd_sc_hd__and3_1
XFILLER_97_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13003_ _12997_/C _12998_/C _13000_/Y _13001_/X vssd1 vssd1 vccd1 vccd1 _13004_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10215_ _10215_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10217_/A sky130_fd_sc_hd__or2_1
X_11195_ _15938_/Q _11197_/C _11023_/X vssd1 vssd1 vccd1 vccd1 _11195_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10146_ _10146_/A vssd1 vssd1 vccd1 vccd1 _15763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16656__61 vssd1 vssd1 vccd1 vccd1 _16656__61/HI _16732_/A sky130_fd_sc_hd__conb_1
XFILLER_121_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10077_ _10179_/A _10077_/B _10081_/A vssd1 vssd1 vccd1 vccd1 _15751_/D sky130_fd_sc_hd__nor3_1
X_14954_ _14954_/A vssd1 vssd1 vccd1 vccd1 _14954_/X sky130_fd_sc_hd__clkbuf_2
X_13905_ _16322_/Q _13908_/C _13853_/X vssd1 vssd1 vccd1 vccd1 _13905_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14885_ _14909_/A _14885_/B _14889_/B vssd1 vssd1 vccd1 vccd1 _16466_/D sky130_fd_sc_hd__nor3_1
X_13836_ _13856_/C vssd1 vssd1 vccd1 vccd1 _13869_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16555_ _16533_/Q _16555_/D vssd1 vssd1 vccd1 vccd1 _16555_/Q sky130_fd_sc_hd__dfxtp_4
X_10979_ _10975_/Y _10976_/X _10978_/Y _10973_/C vssd1 vssd1 vccd1 vccd1 _10981_/B
+ sky130_fd_sc_hd__o211ai_1
X_13767_ _13767_/A _13767_/B vssd1 vssd1 vccd1 vccd1 _13768_/B sky130_fd_sc_hd__nor2_1
X_15506_ _16551_/CLK _15506_/D vssd1 vssd1 vccd1 vccd1 _15506_/Q sky130_fd_sc_hd__dfxtp_1
X_12718_ _16153_/Q _12770_/B _12718_/C vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__and3_1
XFILLER_31_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16486_ _16607_/CLK _16486_/D vssd1 vssd1 vccd1 vccd1 _16486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13698_ _13979_/A vssd1 vssd1 vccd1 vccd1 _13698_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15437_ _16333_/Q _16332_/Q _16331_/Q _15434_/X vssd1 vssd1 vccd1 vccd1 _16612_/D
+ sky130_fd_sc_hd__o31a_1
X_12649_ _12685_/C vssd1 vssd1 vccd1 vccd1 _12692_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15368_ _15884_/Q _15883_/Q _15882_/Q _15363_/X vssd1 vssd1 vccd1 vccd1 _16556_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_144_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14319_ _14316_/Y _14325_/A _14318_/Y _14314_/C vssd1 vssd1 vccd1 vccd1 _14321_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15299_ _15299_/A _15299_/B vssd1 vssd1 vccd1 vccd1 _15300_/A sky130_fd_sc_hd__and2_1
XFILLER_132_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09860_ _15723_/Q vssd1 vssd1 vccd1 vccd1 _09864_/C sky130_fd_sc_hd__inv_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _08811_/A vssd1 vssd1 vccd1 vccd1 _15491_/D sky130_fd_sc_hd__clkbuf_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _09749_/X _09788_/B _09790_/Y vssd1 vssd1 vccd1 vccd1 _15694_/D sky130_fd_sc_hd__o21a_1
XFILLER_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _08630_/X _08733_/B _08736_/B _08741_/Y vssd1 vssd1 vccd1 vccd1 _15476_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08673_ _10833_/B vssd1 vssd1 vccd1 vccd1 _10285_/C sky130_fd_sc_hd__buf_6
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09225_ _15586_/Q _09231_/C _09063_/X vssd1 vssd1 vccd1 vccd1 _09225_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09156_ _10112_/A vssd1 vssd1 vccd1 vccd1 _10065_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08107_ _08108_/A _16703_/A _15282_/C vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__o21a_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09087_ _10276_/A vssd1 vssd1 vccd1 vccd1 _09087_/X sky130_fd_sc_hd__clkbuf_2
X_08038_ _08038_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _08039_/B sky130_fd_sc_hd__nand2_1
XFILLER_123_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10000_ _09994_/C _09995_/C _09997_/Y _10004_/A vssd1 vssd1 vccd1 vccd1 _10004_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_67_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09989_ _10430_/A vssd1 vssd1 vccd1 vccd1 _10340_/A sky130_fd_sc_hd__buf_2
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11951_ _11951_/A _11960_/B vssd1 vssd1 vccd1 vccd1 _11954_/A sky130_fd_sc_hd__or2_1
XFILLER_85_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10902_ _10902_/A _10902_/B _10902_/C vssd1 vssd1 vccd1 vccd1 _10903_/C sky130_fd_sc_hd__nand3_1
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11882_ _11882_/A vssd1 vssd1 vccd1 vccd1 _16033_/D sky130_fd_sc_hd__clkbuf_1
X_14670_ _14671_/B _14671_/C _14669_/X vssd1 vssd1 vccd1 vccd1 _14672_/B sky130_fd_sc_hd__o21ai_1
XFILLER_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13621_ _13621_/A vssd1 vssd1 vccd1 vccd1 _16280_/D sky130_fd_sc_hd__clkbuf_1
X_10833_ _15887_/Q _10833_/B _10844_/C vssd1 vssd1 vccd1 vccd1 _10838_/A sky130_fd_sc_hd__and3_1
XFILLER_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater14 _16554_/Q vssd1 vssd1 vccd1 vccd1 _16118_/CLK sky130_fd_sc_hd__buf_12
X_16340_ _16346_/CLK _16340_/D vssd1 vssd1 vccd1 vccd1 _16340_/Q sky130_fd_sc_hd__dfxtp_1
X_13552_ _13565_/C vssd1 vssd1 vccd1 vccd1 _13573_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10764_ _09308_/X _10762_/B _10716_/X vssd1 vssd1 vccd1 vccd1 _10764_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12503_ _12500_/Y _12501_/X _12502_/Y _12498_/C vssd1 vssd1 vccd1 vccd1 _12505_/B
+ sky130_fd_sc_hd__o211ai_1
X_16271_ _16533_/Q _16271_/D vssd1 vssd1 vccd1 vccd1 _16271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13483_ _13596_/A _13488_/C vssd1 vssd1 vccd1 vccd1 _13483_/X sky130_fd_sc_hd__or2_1
X_10695_ _10738_/A _10695_/B _10695_/C vssd1 vssd1 vccd1 vccd1 _10696_/A sky130_fd_sc_hd__and3_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15222_ _15223_/B _15223_/C _09207_/A vssd1 vssd1 vccd1 vccd1 _15224_/B sky130_fd_sc_hd__o21ai_1
X_12434_ _16113_/Q _12443_/C _12323_/X vssd1 vssd1 vccd1 vccd1 _12434_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15153_ _15153_/A vssd1 vssd1 vccd1 vccd1 _16510_/D sky130_fd_sc_hd__clkbuf_1
X_12365_ _12380_/C vssd1 vssd1 vccd1 vccd1 _12387_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11316_ _15954_/Q _11488_/B _11322_/C vssd1 vssd1 vccd1 vccd1 _11316_/Y sky130_fd_sc_hd__nand3_1
X_14104_ _14104_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14110_/C sky130_fd_sc_hd__nor2_1
XFILLER_99_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15084_ _15082_/Y _15083_/X _15079_/C _15080_/C vssd1 vssd1 vccd1 vccd1 _15086_/B
+ sky130_fd_sc_hd__o211ai_1
X_12296_ _16093_/Q _12516_/B _12296_/C vssd1 vssd1 vccd1 vccd1 _12304_/B sky130_fd_sc_hd__and3_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14035_ _14035_/A _14035_/B _14035_/C vssd1 vssd1 vccd1 vccd1 _14036_/A sky130_fd_sc_hd__and3_1
X_11247_ _11245_/Y _11246_/X _11242_/C _11243_/C vssd1 vssd1 vccd1 vccd1 _11249_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11178_ _12312_/A vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_68_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ _10129_/A _10129_/B _10129_/C vssd1 vssd1 vccd1 vccd1 _10130_/C sky130_fd_sc_hd__nand3_1
X_15986_ _16005_/CLK _15986_/D vssd1 vssd1 vccd1 vccd1 _15986_/Q sky130_fd_sc_hd__dfxtp_1
X_14937_ _14937_/A vssd1 vssd1 vccd1 vccd1 _16474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14868_ _14865_/Y _14866_/X _14867_/Y _14863_/C vssd1 vssd1 vccd1 vccd1 _14870_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16607_ _16607_/CLK _16607_/D vssd1 vssd1 vccd1 vccd1 _16607_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13819_ _13817_/Y _13811_/C _13814_/Y _13824_/A vssd1 vssd1 vccd1 vccd1 _13824_/B
+ sky130_fd_sc_hd__a211oi_1
X_14799_ _14799_/A vssd1 vssd1 vccd1 vccd1 _15027_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16538_ _16570_/CLK _16538_/D vssd1 vssd1 vccd1 vccd1 _16707_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_148_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16469_ _16607_/CLK _16469_/D vssd1 vssd1 vccd1 vccd1 _16469_/Q sky130_fd_sc_hd__dfxtp_1
X_09010_ _09016_/C vssd1 vssd1 vccd1 vccd1 _09028_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09912_ _09912_/A vssd1 vssd1 vccd1 vccd1 _15716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _12849_/A vssd1 vssd1 vccd1 vccd1 _11150_/A sky130_fd_sc_hd__buf_4
XFILLER_140_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _15694_/Q _09781_/C _09683_/X vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__a21oi_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08725_ _08725_/A vssd1 vssd1 vccd1 vccd1 _15473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _08656_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _15460_/D sky130_fd_sc_hd__nor2_1
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08587_ _15235_/B vssd1 vssd1 vccd1 vccd1 _10183_/A sky130_fd_sc_hd__buf_4
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09208_ _09207_/X _09206_/A _09129_/X vssd1 vssd1 vccd1 vccd1 _09208_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10480_ _10494_/C vssd1 vssd1 vccd1 vccd1 _10509_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09139_ _15567_/Q _09220_/B _09139_/C vssd1 vssd1 vccd1 vccd1 _09141_/C sky130_fd_sc_hd__nand3_1
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12150_ _12150_/A vssd1 vssd1 vccd1 vccd1 _16071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11101_ _11101_/A _11101_/B vssd1 vssd1 vccd1 vccd1 _11103_/B sky130_fd_sc_hd__nor2_1
XFILLER_150_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12081_/X sky130_fd_sc_hd__clkbuf_2
X_11032_ _15915_/Q _11084_/B _11039_/C vssd1 vssd1 vccd1 vccd1 _11032_/X sky130_fd_sc_hd__and3_1
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15840_ _16551_/CLK _15840_/D vssd1 vssd1 vccd1 vccd1 _15840_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16626__31 vssd1 vssd1 vccd1 vccd1 _16626__31/HI _16692_/A sky130_fd_sc_hd__conb_1
XFILLER_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15771_ _15791_/CLK _15771_/D vssd1 vssd1 vccd1 vccd1 _15771_/Q sky130_fd_sc_hd__dfxtp_1
X_12983_ _12984_/B _12984_/C _12982_/X vssd1 vssd1 vccd1 vccd1 _12985_/B sky130_fd_sc_hd__o21ai_1
XFILLER_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14722_ _14722_/A vssd1 vssd1 vccd1 vccd1 _14760_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11934_ _11934_/A vssd1 vssd1 vccd1 vccd1 _16041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14653_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14768_/A sky130_fd_sc_hd__clkbuf_2
X_11865_ _11865_/A _11865_/B _11865_/C vssd1 vssd1 vccd1 vccd1 _11866_/C sky130_fd_sc_hd__nand3_1
XFILLER_26_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13604_ _13617_/C vssd1 vssd1 vccd1 vccd1 _13625_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10816_ _10816_/A _10816_/B vssd1 vssd1 vccd1 vccd1 _10823_/C sky130_fd_sc_hd__nor2_1
XFILLER_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11796_ _11832_/A _11796_/B _11796_/C vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__and3_1
X_14584_ _14581_/Y _14582_/X _14583_/Y _14579_/C vssd1 vssd1 vccd1 vccd1 _14586_/B
+ sky130_fd_sc_hd__o211ai_1
X_16323_ _16346_/CLK _16323_/D vssd1 vssd1 vccd1 vccd1 _16323_/Q sky130_fd_sc_hd__dfxtp_1
X_13535_ _13533_/Y _13526_/C _13530_/Y _13540_/A vssd1 vssd1 vccd1 vccd1 _13540_/B
+ sky130_fd_sc_hd__a211oi_1
X_10747_ _10747_/A vssd1 vssd1 vccd1 vccd1 _15871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16254_ _16261_/CLK _16254_/D vssd1 vssd1 vccd1 vccd1 _16254_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10678_ _15862_/Q _10685_/C _09629_/A vssd1 vssd1 vccd1 vccd1 _10681_/B sky130_fd_sc_hd__a21o_1
X_13466_ _16259_/Q _13631_/B _13473_/C vssd1 vssd1 vccd1 vccd1 _13466_/X sky130_fd_sc_hd__and3_1
XFILLER_145_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15205_ _15205_/A _15205_/B _15205_/C vssd1 vssd1 vccd1 vccd1 _15206_/A sky130_fd_sc_hd__and3_1
X_12417_ _12418_/B _12418_/C _12416_/X vssd1 vssd1 vccd1 vccd1 _12419_/B sky130_fd_sc_hd__o21ai_1
X_16185_ _16555_/Q _16185_/D vssd1 vssd1 vccd1 vccd1 _16185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13397_ _13397_/A vssd1 vssd1 vccd1 vccd1 _16248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15136_ _15134_/Y _15135_/X _15131_/C _15132_/C vssd1 vssd1 vccd1 vccd1 _15138_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_127_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12348_ _12345_/Y _12354_/A _12347_/Y _12343_/C vssd1 vssd1 vccd1 vccd1 _12350_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15067_ _16486_/Q _16485_/Q _16484_/Q _14900_/X vssd1 vssd1 vccd1 vccd1 _16496_/D
+ sky130_fd_sc_hd__o31a_1
X_12279_ _16091_/Q _12501_/B _12287_/C vssd1 vssd1 vccd1 vccd1 _12279_/X sky130_fd_sc_hd__and3_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14018_ _14016_/Y _14017_/X _14012_/C _14013_/C vssd1 vssd1 vccd1 vccd1 _14020_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15969_ _16005_/CLK _15969_/D vssd1 vssd1 vccd1 vccd1 _15969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08510_ _08542_/A _08510_/B vssd1 vssd1 vccd1 vccd1 _08537_/B sky130_fd_sc_hd__nor2_2
X_09490_ _15623_/Q _15622_/Q _15621_/Q _09314_/X vssd1 vssd1 vccd1 vccd1 _15633_/D
+ sky130_fd_sc_hd__o31a_1
X_08441_ _08441_/A _08441_/B vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08372_ _08372_/A _08372_/B vssd1 vssd1 vccd1 vccd1 _08454_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09826_ _15702_/Q _10300_/C _09836_/C vssd1 vssd1 vccd1 vccd1 _09826_/X sky130_fd_sc_hd__and3_1
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09757_ _15677_/Q _15676_/Q _15675_/Q _09756_/X vssd1 vssd1 vccd1 vccd1 _15687_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _15338_/A vssd1 vssd1 vccd1 vccd1 _08708_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09688_/A _09688_/B vssd1 vssd1 vccd1 vccd1 _09688_/X sky130_fd_sc_hd__or2_1
XFILLER_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _10755_/B vssd1 vssd1 vccd1 vccd1 _09699_/A sky130_fd_sc_hd__buf_2
XFILLER_70_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11648_/Y _11641_/C _11643_/Y _11644_/X vssd1 vssd1 vccd1 vccd1 _11651_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ _10598_/Y _10599_/X _10600_/Y _10596_/C vssd1 vssd1 vccd1 vccd1 _10603_/B
+ sky130_fd_sc_hd__o211ai_1
X_11581_ _11582_/B _11582_/C _11582_/A vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__a21o_1
XFILLER_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10532_ _10546_/C vssd1 vssd1 vccd1 vccd1 _10559_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13320_ _13354_/A _13320_/B _13320_/C vssd1 vssd1 vccd1 vccd1 _13321_/A sky130_fd_sc_hd__and3_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10463_ _15821_/Q _10463_/B _10463_/C vssd1 vssd1 vccd1 vccd1 _10464_/B sky130_fd_sc_hd__and3_1
X_13251_ _14095_/A vssd1 vssd1 vccd1 vccd1 _13474_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ _12202_/A vssd1 vssd1 vccd1 vccd1 _16079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13182_ _13182_/A vssd1 vssd1 vccd1 vccd1 _16217_/D sky130_fd_sc_hd__clkbuf_1
X_10394_ _15810_/Q _10402_/C _10393_/X vssd1 vssd1 vccd1 vccd1 _10394_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12133_ _13264_/A vssd1 vssd1 vccd1 vccd1 _12133_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12064_ _16061_/Q _12065_/C _12007_/X vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__a21oi_1
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11015_ _11036_/A _11015_/B _11015_/C vssd1 vssd1 vccd1 vccd1 _11016_/A sky130_fd_sc_hd__and3_1
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15823_ _16595_/CLK _15823_/D vssd1 vssd1 vccd1 vccd1 _15823_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15754_ _15791_/CLK _15754_/D vssd1 vssd1 vccd1 vccd1 _15754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12966_ _16188_/Q _12975_/C _12850_/X vssd1 vssd1 vccd1 vccd1 _12966_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14705_ _14702_/Y _14703_/X _14704_/Y _14700_/C vssd1 vssd1 vccd1 vccd1 _14707_/B
+ sky130_fd_sc_hd__o211ai_1
X_11917_ _11918_/B _11918_/C _11918_/A vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__a21o_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _15791_/CLK _15685_/D vssd1 vssd1 vccd1 vccd1 _15685_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12894_/Y _12895_/X _12896_/Y _12892_/C vssd1 vssd1 vccd1 vccd1 _12899_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14636_ _14651_/A _14636_/B _14636_/C vssd1 vssd1 vccd1 vccd1 _14637_/A sky130_fd_sc_hd__and3_1
X_11848_ _11846_/A _11846_/B _11847_/X vssd1 vssd1 vccd1 vccd1 _16028_/D sky130_fd_sc_hd__a21oi_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14567_ _14851_/A vssd1 vssd1 vccd1 vccd1 _14567_/X sky130_fd_sc_hd__clkbuf_4
X_11779_ _16020_/Q _11891_/B _11779_/C vssd1 vssd1 vccd1 vccd1 _11787_/A sky130_fd_sc_hd__and3_1
XFILLER_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16306_ _16346_/CLK _16306_/D vssd1 vssd1 vccd1 vccd1 _16306_/Q sky130_fd_sc_hd__dfxtp_1
X_13518_ _13518_/A vssd1 vssd1 vccd1 vccd1 _16265_/D sky130_fd_sc_hd__clkbuf_1
X_14498_ _14498_/A vssd1 vssd1 vccd1 vccd1 _16405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16237_ _16237_/CLK _16237_/D vssd1 vssd1 vccd1 vccd1 _16237_/Q sky130_fd_sc_hd__dfxtp_1
X_13449_ _13449_/A vssd1 vssd1 vccd1 vccd1 _16255_/D sky130_fd_sc_hd__clkbuf_1
X_16168_ _16237_/CLK _16168_/D vssd1 vssd1 vccd1 vccd1 _16168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15119_ _15119_/A vssd1 vssd1 vccd1 vccd1 _16504_/D sky130_fd_sc_hd__clkbuf_1
X_08990_ _15533_/Q _08991_/C _08989_/X vssd1 vssd1 vccd1 vccd1 _08992_/A sky130_fd_sc_hd__a21oi_1
X_16099_ _16118_/CLK _16099_/D vssd1 vssd1 vccd1 vccd1 _16099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07941_ _07941_/A _07941_/B vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07872_ _07872_/A _07872_/B vssd1 vssd1 vccd1 vccd1 _07873_/B sky130_fd_sc_hd__nand2_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09611_ _09656_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _09611_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09542_ _09595_/A _09542_/B _09546_/A vssd1 vssd1 vccd1 vccd1 _15643_/D sky130_fd_sc_hd__nor3_1
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09473_ _15632_/Q _09472_/C _09383_/X vssd1 vssd1 vccd1 vccd1 _09474_/B sky130_fd_sc_hd__a21o_1
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08424_ input8/X vssd1 vssd1 vccd1 vccd1 _08526_/A sky130_fd_sc_hd__inv_2
XFILLER_12_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08355_ _08355_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08359_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08286_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08287_/B sky130_fd_sc_hd__xor2_1
XFILLER_137_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09809_ _09809_/A _09809_/B _09809_/C vssd1 vssd1 vccd1 vccd1 _09810_/C sky130_fd_sc_hd__nand3_1
XFILLER_74_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12820_ _16168_/Q _12828_/C _12598_/X vssd1 vssd1 vccd1 vccd1 _12823_/B sky130_fd_sc_hd__a21o_1
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12751_/A vssd1 vssd1 vccd1 vccd1 _12788_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11702_/A vssd1 vssd1 vccd1 vccd1 _16008_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15470_ _16551_/CLK _15470_/D vssd1 vssd1 vccd1 vccd1 _15470_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12682_/A vssd1 vssd1 vccd1 vccd1 _16146_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14421_ _16394_/Q _14591_/B _14427_/C vssd1 vssd1 vccd1 vccd1 _14421_/Y sky130_fd_sc_hd__nand3_1
X_11633_ _11634_/B _11634_/C _11634_/A vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__a21o_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14352_ _14350_/Y _14351_/X _14347_/C _14348_/C vssd1 vssd1 vccd1 vccd1 _14354_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ _11617_/A _11569_/C vssd1 vssd1 vccd1 vccd1 _11564_/X sky130_fd_sc_hd__or2_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _13303_/A vssd1 vssd1 vccd1 vccd1 _16234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10515_ _15830_/Q _10517_/C _10360_/X vssd1 vssd1 vccd1 vccd1 _10518_/A sky130_fd_sc_hd__a21oi_1
X_11495_ _15979_/Q _11495_/B _11500_/C vssd1 vssd1 vccd1 vccd1 _11495_/Y sky130_fd_sc_hd__nand3_1
X_14283_ _16375_/Q _14323_/C _14060_/X vssd1 vssd1 vccd1 vccd1 _14286_/B sky130_fd_sc_hd__a21oi_1
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16022_ _16118_/CLK _16022_/D vssd1 vssd1 vccd1 vccd1 _16022_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10446_ _15819_/Q _10446_/B _10457_/C vssd1 vssd1 vccd1 vccd1 _10446_/X sky130_fd_sc_hd__and3_1
X_13234_ _16226_/Q _13342_/B _13235_/C vssd1 vssd1 vccd1 vccd1 _13234_/X sky130_fd_sc_hd__and3_1
XFILLER_108_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _13166_/B _13166_/C _13166_/A vssd1 vssd1 vccd1 vccd1 _13167_/B sky130_fd_sc_hd__a21o_1
X_10377_ _10402_/C vssd1 vssd1 vccd1 vccd1 _10408_/C sky130_fd_sc_hd__clkbuf_2
X_12116_ _12683_/A vssd1 vssd1 vccd1 vccd1 _12230_/A sky130_fd_sc_hd__buf_2
XFILLER_123_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13096_ _13377_/A vssd1 vssd1 vccd1 vccd1 _13219_/A sky130_fd_sc_hd__buf_2
XFILLER_78_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12047_ _12045_/Y _12041_/C _12043_/Y _12044_/X vssd1 vssd1 vccd1 vccd1 _12048_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15806_ _16595_/CLK _15806_/D vssd1 vssd1 vccd1 vccd1 _15806_/Q sky130_fd_sc_hd__dfxtp_2
X_13998_ _14035_/A _13998_/B _13998_/C vssd1 vssd1 vccd1 vccd1 _13999_/A sky130_fd_sc_hd__and3_1
X_15737_ _16551_/CLK _15737_/D vssd1 vssd1 vccd1 vccd1 _15737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ _12949_/A vssd1 vssd1 vccd1 vccd1 _16184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15668_ _15791_/CLK _15668_/D vssd1 vssd1 vccd1 vccd1 _15668_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14619_ _14640_/C vssd1 vssd1 vccd1 vccd1 _14655_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15599_ _16570_/CLK _15599_/D vssd1 vssd1 vccd1 vccd1 _15599_/Q sky130_fd_sc_hd__dfxtp_2
X_08140_ _09905_/C _08140_/B vssd1 vssd1 vccd1 vccd1 _08140_/X sky130_fd_sc_hd__or2_1
X_08071_ _16505_/Q vssd1 vssd1 vccd1 vccd1 _15013_/A sky130_fd_sc_hd__clkinv_2
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08973_ _15530_/Q _09053_/B _08978_/C vssd1 vssd1 vccd1 vccd1 _08980_/A sky130_fd_sc_hd__and3_1
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07924_ _16603_/Q vssd1 vssd1 vccd1 vccd1 _13435_/A sky130_fd_sc_hd__clkinv_2
XFILLER_96_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07855_ _07855_/A vssd1 vssd1 vccd1 vccd1 _08678_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_83_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07786_ _07787_/A vssd1 vssd1 vccd1 vccd1 _07786_/Y sky130_fd_sc_hd__inv_2
X_09525_ _09517_/Y _09519_/X _09521_/B vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__o21a_1
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09456_ _15630_/Q _09458_/C _09369_/X vssd1 vssd1 vccd1 vccd1 _09456_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _08407_/A _08407_/B vssd1 vssd1 vccd1 vccd1 _08410_/A sky130_fd_sc_hd__xnor2_1
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09387_ _09381_/Y _09385_/X _09386_/Y vssd1 vssd1 vccd1 vccd1 _15611_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ _08338_/A _08338_/B vssd1 vssd1 vccd1 vccd1 _08440_/A sky130_fd_sc_hd__xor2_4
XFILLER_137_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08269_ _08386_/A _08386_/B vssd1 vssd1 vccd1 vccd1 _08273_/A sky130_fd_sc_hd__xnor2_1
XFILLER_138_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10300_ _15792_/Q _10307_/B _10300_/C vssd1 vssd1 vccd1 vccd1 _10300_/X sky130_fd_sc_hd__and3_1
X_11280_ _11278_/A _11278_/B _11279_/X vssd1 vssd1 vccd1 vccd1 _15948_/D sky130_fd_sc_hd__a21oi_1
XFILLER_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10231_ _10247_/C vssd1 vssd1 vccd1 vccd1 _10261_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10162_ _10271_/A _10162_/B vssd1 vssd1 vccd1 vccd1 _10162_/X sky130_fd_sc_hd__or2_1
XFILLER_121_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10093_ _15755_/Q _10301_/C _10099_/C vssd1 vssd1 vccd1 vccd1 _10093_/Y sky130_fd_sc_hd__nand3_1
XFILLER_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14970_ _14970_/A _14970_/B _14970_/C vssd1 vssd1 vccd1 vccd1 _14971_/C sky130_fd_sc_hd__nand3_1
XFILLER_94_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13921_ input5/X vssd1 vssd1 vccd1 vccd1 _15048_/A sky130_fd_sc_hd__buf_4
X_13852_ _13852_/A vssd1 vssd1 vccd1 vccd1 _16312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ _13032_/A _12808_/C vssd1 vssd1 vccd1 vccd1 _12803_/X sky130_fd_sc_hd__or2_1
X_16571_ _16595_/CLK _16571_/D vssd1 vssd1 vccd1 vccd1 _16571_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13783_ _16303_/Q _13948_/B _13793_/C vssd1 vssd1 vccd1 vccd1 _13789_/A sky130_fd_sc_hd__and3_1
X_10995_ _10995_/A _10995_/B vssd1 vssd1 vccd1 vccd1 _11001_/C sky130_fd_sc_hd__nor2_1
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15522_ _16551_/CLK _15522_/D vssd1 vssd1 vccd1 vccd1 _15522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12734_ _12731_/Y _12732_/X _12733_/Y _12729_/C vssd1 vssd1 vccd1 vccd1 _12736_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _16570_/CLK _15453_/D vssd1 vssd1 vccd1 vccd1 _15453_/Q sky130_fd_sc_hd__dfxtp_1
X_12665_ _12659_/C _12660_/C _12662_/Y _12663_/X vssd1 vssd1 vccd1 vccd1 _12666_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14404_ _14404_/A vssd1 vssd1 vccd1 vccd1 _16391_/D sky130_fd_sc_hd__clkbuf_1
X_11616_ _11616_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11621_/C sky130_fd_sc_hd__nor2_1
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15384_ _15415_/A vssd1 vssd1 vccd1 vccd1 _15409_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12596_ _16135_/Q _12818_/B _12607_/C vssd1 vssd1 vccd1 vccd1 _12602_/A sky130_fd_sc_hd__and3_1
X_14335_ _14335_/A vssd1 vssd1 vccd1 vccd1 _14351_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11547_ _11547_/A _11547_/B _11547_/C vssd1 vssd1 vccd1 vccd1 _11548_/A sky130_fd_sc_hd__and3_1
XFILLER_144_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14266_ _16373_/Q _14268_/C _14265_/X vssd1 vssd1 vccd1 vccd1 _14269_/A sky130_fd_sc_hd__a21oi_1
X_11478_ _15978_/Q _11480_/C _11306_/X vssd1 vssd1 vccd1 vccd1 _11478_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16005_ _16005_/CLK _16005_/D vssd1 vssd1 vccd1 vccd1 _16005_/Q sky130_fd_sc_hd__dfxtp_1
X_13217_ _16223_/Q _13257_/C _13216_/X vssd1 vssd1 vccd1 vccd1 _13219_/B sky130_fd_sc_hd__a21oi_1
X_10429_ _10429_/A _10429_/B _10436_/A vssd1 vssd1 vccd1 vccd1 _15814_/D sky130_fd_sc_hd__nor3_1
XFILLER_124_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14197_ _14197_/A _14197_/B _14197_/C vssd1 vssd1 vccd1 vccd1 _14198_/A sky130_fd_sc_hd__and3_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _13146_/A _13146_/B _13147_/X vssd1 vssd1 vccd1 vccd1 _16212_/D sky130_fd_sc_hd__a21oi_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13079_ _13077_/Y _13072_/C _13074_/Y _13084_/A vssd1 vssd1 vccd1 vccd1 _13084_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_112_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09310_ _14895_/A vssd1 vssd1 vccd1 vccd1 _11850_/A sky130_fd_sc_hd__buf_6
XFILLER_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ _15358_/A vssd1 vssd1 vccd1 vccd1 _09744_/A sky130_fd_sc_hd__buf_2
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09172_ _09178_/C vssd1 vssd1 vccd1 vccd1 _09192_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_08123_ _07949_/A _07949_/B _07948_/A vssd1 vssd1 vccd1 vccd1 _08138_/A sky130_fd_sc_hd__o21a_1
XFILLER_135_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ _16590_/Q vssd1 vssd1 vccd1 vccd1 _12704_/A sky130_fd_sc_hd__clkinv_2
XFILLER_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08956_ _09119_/A _08963_/C vssd1 vssd1 vccd1 vccd1 _08956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07907_ _16612_/Q vssd1 vssd1 vccd1 vccd1 _13943_/A sky130_fd_sc_hd__clkinv_4
X_08887_ _09756_/A vssd1 vssd1 vccd1 vccd1 _08887_/X sky130_fd_sc_hd__buf_2
XFILLER_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07838_ _07842_/A vssd1 vssd1 vccd1 vccd1 _07838_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07769_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07774_/A sky130_fd_sc_hd__buf_12
X_09508_ _09506_/Y _09513_/A _09501_/C _09502_/C vssd1 vssd1 vccd1 vccd1 _09510_/B
+ sky130_fd_sc_hd__o211a_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ _14858_/A vssd1 vssd1 vccd1 vccd1 _15034_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09438_/X _09436_/B _09431_/X vssd1 vssd1 vccd1 vccd1 _09439_/Y sky130_fd_sc_hd__a21oi_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _16114_/Q _12622_/B _12456_/C vssd1 vssd1 vccd1 vccd1 _12450_/Y sky130_fd_sc_hd__nand3_1
XFILLER_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _15967_/Q _11444_/C _11233_/X vssd1 vssd1 vccd1 vccd1 _11403_/B sky130_fd_sc_hd__a21oi_1
X_12381_ _12379_/Y _12380_/X _12376_/C _12377_/C vssd1 vssd1 vccd1 vccd1 _12383_/B
+ sky130_fd_sc_hd__o211ai_1
X_14120_ _16352_/Q _14127_/C _14008_/X vssd1 vssd1 vccd1 vccd1 _14123_/B sky130_fd_sc_hd__a21o_1
X_11332_ _11332_/A _11336_/C vssd1 vssd1 vccd1 vccd1 _11332_/X sky130_fd_sc_hd__or2_1
XFILLER_125_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ _14053_/B _14053_/C _13829_/X vssd1 vssd1 vccd1 vccd1 _14054_/B sky130_fd_sc_hd__o21ai_1
X_11263_ _11261_/Y _11256_/C _11258_/Y _11259_/X vssd1 vssd1 vccd1 vccd1 _11264_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_106_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _13000_/Y _13001_/X _12997_/C _12998_/C vssd1 vssd1 vccd1 vccd1 _13004_/B
+ sky130_fd_sc_hd__o211ai_1
X_10214_ _15776_/Q _10463_/B _10214_/C vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__and3_1
X_11194_ _11194_/A vssd1 vssd1 vccd1 vccd1 _15936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10145_ _10145_/A _10145_/B _10145_/C vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__and3_1
XFILLER_97_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10076_ _15753_/Q _10178_/B _10076_/C vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__and3_1
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14953_ _15007_/A vssd1 vssd1 vccd1 vccd1 _14992_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13904_ _13904_/A vssd1 vssd1 vccd1 vccd1 _16320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14884_ _14882_/Y _14878_/C _14880_/Y _14889_/A vssd1 vssd1 vccd1 vccd1 _14889_/B
+ sky130_fd_sc_hd__a211oi_1
X_16671__76 vssd1 vssd1 vccd1 vccd1 _16671__76/HI _16747_/A sky130_fd_sc_hd__conb_1
XFILLER_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13835_ _13848_/C vssd1 vssd1 vccd1 vccd1 _13856_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16554_ _16555_/Q _16554_/D vssd1 vssd1 vccd1 vccd1 _16554_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13766_ _13766_/A _13774_/B vssd1 vssd1 vccd1 vccd1 _13768_/A sky130_fd_sc_hd__or2_1
X_10978_ _15906_/Q _11205_/B _10985_/C vssd1 vssd1 vccd1 vccd1 _10978_/Y sky130_fd_sc_hd__nand3_1
XFILLER_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _16551_/CLK _15505_/D vssd1 vssd1 vccd1 vccd1 _15505_/Q sky130_fd_sc_hd__dfxtp_1
X_12717_ _16153_/Q _12726_/C _12605_/X vssd1 vssd1 vccd1 vccd1 _12717_/Y sky130_fd_sc_hd__a21oi_1
X_16485_ _16607_/CLK _16485_/D vssd1 vssd1 vccd1 vccd1 _16485_/Q sky130_fd_sc_hd__dfxtp_1
X_13697_ _13697_/A vssd1 vssd1 vccd1 vccd1 _16290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15436_ _16325_/Q _16324_/Q _16323_/Q _15434_/X vssd1 vssd1 vccd1 vccd1 _16611_/D
+ sky130_fd_sc_hd__o31a_1
X_12648_ _12670_/C vssd1 vssd1 vccd1 vccd1 _12685_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15367_ _16555_/Q _15367_/B vssd1 vssd1 vccd1 vccd1 _16555_/D sky130_fd_sc_hd__nor2_1
X_12579_ _12579_/A _12586_/B vssd1 vssd1 vccd1 vccd1 _12581_/A sky130_fd_sc_hd__or2_1
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14318_ _16379_/Q _14318_/B _14323_/C vssd1 vssd1 vccd1 vccd1 _14318_/Y sky130_fd_sc_hd__nand3_1
X_15298_ _15299_/A _15299_/B vssd1 vssd1 vccd1 vccd1 _15301_/A sky130_fd_sc_hd__or2_1
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14249_ _14249_/A vssd1 vssd1 vccd1 vccd1 _16369_/D sky130_fd_sc_hd__clkbuf_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08810_ _08940_/A _08810_/B _08810_/C vssd1 vssd1 vccd1 vccd1 _08811_/A sky130_fd_sc_hd__and3_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09658_/X _09788_/B _09750_/X vssd1 vssd1 vccd1 vccd1 _09790_/Y sky130_fd_sc_hd__a21oi_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08741_ _08916_/A _08752_/C vssd1 vssd1 vccd1 vccd1 _08741_/Y sky130_fd_sc_hd__nor2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08672_ _14848_/A vssd1 vssd1 vccd1 vccd1 _10833_/B sky130_fd_sc_hd__buf_2
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _09224_/A vssd1 vssd1 vccd1 vccd1 _15581_/D sky130_fd_sc_hd__clkbuf_1
X_09155_ _09153_/A _09153_/B _09154_/X vssd1 vssd1 vccd1 vccd1 _15565_/D sky130_fd_sc_hd__a21oi_1
XFILLER_148_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08106_ _08678_/C _08106_/B vssd1 vssd1 vccd1 vccd1 _15282_/C sky130_fd_sc_hd__xnor2_2
X_09086_ _09086_/A _09086_/B vssd1 vssd1 vccd1 vccd1 _15550_/D sky130_fd_sc_hd__nor2_1
XFILLER_135_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08037_ _08038_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _08039_/A sky130_fd_sc_hd__or2_1
XFILLER_150_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09988_ _10055_/A _09988_/B _09994_/A vssd1 vssd1 vccd1 vccd1 _15733_/D sky130_fd_sc_hd__nor3_1
XFILLER_88_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08939_ _08939_/A _08939_/B _08939_/C vssd1 vssd1 vccd1 vccd1 _08940_/C sky130_fd_sc_hd__nand3_1
XFILLER_45_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11950_ _16045_/Q _11950_/B _11950_/C vssd1 vssd1 vccd1 vccd1 _11960_/B sky130_fd_sc_hd__and3_1
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10901_ _10902_/B _10902_/C _10902_/A vssd1 vssd1 vccd1 vccd1 _10903_/B sky130_fd_sc_hd__a21o_1
XFILLER_123_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11881_ _11888_/A _11881_/B _11881_/C vssd1 vssd1 vccd1 vccd1 _11882_/A sky130_fd_sc_hd__and3_1
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ _13635_/A _13620_/B _13620_/C vssd1 vssd1 vccd1 vccd1 _13621_/A sky130_fd_sc_hd__and3_1
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10832_ _15887_/Q _10878_/C _10673_/X vssd1 vssd1 vccd1 vccd1 _10834_/B sky130_fd_sc_hd__a21oi_1
XFILLER_53_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater15 _16555_/Q vssd1 vssd1 vccd1 vccd1 _16237_/CLK sky130_fd_sc_hd__buf_12
X_13551_ _13551_/A vssd1 vssd1 vccd1 vccd1 _13565_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10763_ _09301_/X _10756_/B _10759_/B _10762_/Y vssd1 vssd1 vccd1 vccd1 _15874_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_13_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12502_ _16122_/Q _12622_/B _12510_/C vssd1 vssd1 vccd1 vccd1 _12502_/Y sky130_fd_sc_hd__nand3_1
X_16270_ _16533_/Q _16270_/D vssd1 vssd1 vccd1 vccd1 _16270_/Q sky130_fd_sc_hd__dfxtp_2
X_13482_ _13482_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _13488_/C sky130_fd_sc_hd__nor2_1
X_10694_ _10692_/Y _10688_/C _10690_/Y _10691_/X vssd1 vssd1 vccd1 vccd1 _10695_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15221_ _15221_/A vssd1 vssd1 vccd1 vccd1 _15258_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12433_ _12433_/A vssd1 vssd1 vccd1 vccd1 _16111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ _15152_/A _15152_/B _15152_/C vssd1 vssd1 vccd1 vccd1 _15153_/A sky130_fd_sc_hd__and3_1
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12364_ _12364_/A vssd1 vssd1 vccd1 vccd1 _12380_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14103_ _14103_/A _14103_/B vssd1 vssd1 vccd1 vccd1 _14104_/B sky130_fd_sc_hd__nor2_1
X_11315_ _15955_/Q _11367_/B _11322_/C vssd1 vssd1 vccd1 vccd1 _11315_/X sky130_fd_sc_hd__and3_1
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15083_ _16500_/Q _15241_/B _15083_/C vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__and3_1
X_12295_ _13423_/A vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_4_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14034_ _14032_/Y _14027_/C _14030_/Y _14031_/X vssd1 vssd1 vccd1 vccd1 _14035_/C
+ sky130_fd_sc_hd__a211o_1
X_11246_ _15945_/Q _11353_/B _11246_/C vssd1 vssd1 vccd1 vccd1 _11246_/X sky130_fd_sc_hd__and3_1
XFILLER_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ input9/X vssd1 vssd1 vccd1 vccd1 _12312_/A sky130_fd_sc_hd__clkbuf_4
X_10128_ _10129_/B _10129_/C _10129_/A vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__a21o_1
X_15985_ _16005_/CLK _15985_/D vssd1 vssd1 vccd1 vccd1 _15985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10059_ _10059_/A _10059_/B vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__nor2_1
X_14936_ _14936_/A _14936_/B _14936_/C vssd1 vssd1 vccd1 vccd1 _14937_/A sky130_fd_sc_hd__and3_1
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14867_ _16464_/Q _14982_/B _14867_/C vssd1 vssd1 vccd1 vccd1 _14867_/Y sky130_fd_sc_hd__nand3_1
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16606_ _16607_/CLK _16606_/D vssd1 vssd1 vccd1 vccd1 _16606_/Q sky130_fd_sc_hd__dfxtp_1
X_13818_ _13814_/Y _13824_/A _13817_/Y _13811_/C vssd1 vssd1 vccd1 vccd1 _13820_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14798_ _16455_/Q _14808_/C _14574_/X vssd1 vssd1 vccd1 vccd1 _14798_/Y sky130_fd_sc_hd__a21oi_1
X_16537_ _16570_/CLK _16537_/D vssd1 vssd1 vccd1 vccd1 _16706_/A sky130_fd_sc_hd__dfxtp_1
X_13749_ _13749_/A vssd1 vssd1 vccd1 vccd1 _16297_/D sky130_fd_sc_hd__clkbuf_1
X_16468_ _16607_/CLK _16468_/D vssd1 vssd1 vccd1 vccd1 _16468_/Q sky130_fd_sc_hd__dfxtp_1
X_15419_ _16213_/Q _16212_/Q _16211_/Q _15416_/X vssd1 vssd1 vccd1 vccd1 _16597_/D
+ sky130_fd_sc_hd__o31a_1
X_16399_ input11/X _16399_/D vssd1 vssd1 vccd1 vccd1 _16399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09911_ _09951_/A _09911_/B _09911_/C vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__and3_1
XFILLER_104_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09842_ _15704_/Q _09845_/C _09699_/A vssd1 vssd1 vccd1 vccd1 _09846_/A sky130_fd_sc_hd__a21oi_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09841_/A _09773_/B _09776_/B vssd1 vssd1 vccd1 vccd1 _15690_/D sky130_fd_sc_hd__nor3_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08724_ _15304_/A _08724_/B _08724_/C vssd1 vssd1 vccd1 vccd1 _08725_/A sky130_fd_sc_hd__and3_1
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _08654_/X _08646_/A _15312_/A vssd1 vssd1 vccd1 vccd1 _08656_/B sky130_fd_sc_hd__o21ai_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08586_ _12655_/A vssd1 vssd1 vccd1 vccd1 _15235_/B sky130_fd_sc_hd__buf_2
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09207_ _09207_/A vssd1 vssd1 vccd1 vccd1 _09207_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09138_ _15567_/Q _09139_/C _09014_/X vssd1 vssd1 vccd1 vccd1 _09141_/B sky130_fd_sc_hd__a21o_1
XFILLER_136_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09069_ _15551_/Q _09070_/C _08989_/X vssd1 vssd1 vccd1 vccd1 _09071_/A sky130_fd_sc_hd__a21oi_1
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11100_ _11100_/A _11109_/B vssd1 vssd1 vccd1 vccd1 _11103_/A sky130_fd_sc_hd__or2_1
X_12080_ _12118_/C vssd1 vssd1 vccd1 vccd1 _12125_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _15915_/Q _11039_/C _10919_/X vssd1 vssd1 vccd1 vccd1 _11031_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15770_ _15791_/CLK _15770_/D vssd1 vssd1 vccd1 vccd1 _15770_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12982_ _13264_/A vssd1 vssd1 vccd1 vccd1 _12982_/X sky130_fd_sc_hd__buf_2
XFILLER_17_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14721_ _14719_/A _14719_/B _14720_/X vssd1 vssd1 vccd1 vccd1 _16440_/D sky130_fd_sc_hd__a21oi_1
X_11933_ _11940_/A _11933_/B _11933_/C vssd1 vssd1 vccd1 vccd1 _11934_/A sky130_fd_sc_hd__and3_1
XFILLER_73_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16641__46 vssd1 vssd1 vccd1 vccd1 _16641__46/HI _16717_/A sky130_fd_sc_hd__conb_1
XFILLER_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14652_ _14652_/A vssd1 vssd1 vccd1 vccd1 _16429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ _11865_/B _11865_/C _11865_/A vssd1 vssd1 vccd1 vccd1 _11866_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13603_ _13603_/A vssd1 vssd1 vccd1 vccd1 _13617_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10815_ _11384_/A vssd1 vssd1 vccd1 vccd1 _11049_/A sky130_fd_sc_hd__clkbuf_2
X_14583_ _16419_/Q _14697_/B _14583_/C vssd1 vssd1 vccd1 vccd1 _14583_/Y sky130_fd_sc_hd__nand3_1
X_11795_ _12018_/A _11795_/B _11795_/C vssd1 vssd1 vccd1 vccd1 _11796_/C sky130_fd_sc_hd__or3_1
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16322_ _16346_/CLK _16322_/D vssd1 vssd1 vccd1 vccd1 _16322_/Q sky130_fd_sc_hd__dfxtp_1
X_13534_ _13530_/Y _13540_/A _13533_/Y _13526_/C vssd1 vssd1 vccd1 vccd1 _13536_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10746_ _10801_/A _10746_/B _10746_/C vssd1 vssd1 vccd1 vccd1 _10747_/A sky130_fd_sc_hd__and3_1
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16253_ _16261_/CLK _16253_/D vssd1 vssd1 vccd1 vccd1 _16253_/Q sky130_fd_sc_hd__dfxtp_1
X_13465_ _16259_/Q _13473_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13465_/Y sky130_fd_sc_hd__a21oi_1
X_10677_ _10740_/A vssd1 vssd1 vccd1 vccd1 _10738_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ _15202_/Y _15198_/C _15200_/Y _15201_/X vssd1 vssd1 vccd1 vccd1 _15205_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12416_ _13264_/A vssd1 vssd1 vccd1 vccd1 _12416_/X sky130_fd_sc_hd__clkbuf_2
X_16184_ _16237_/CLK _16184_/D vssd1 vssd1 vccd1 vccd1 _16184_/Q sky130_fd_sc_hd__dfxtp_1
X_13396_ _13412_/A _13396_/B _13396_/C vssd1 vssd1 vccd1 vccd1 _13397_/A sky130_fd_sc_hd__and3_1
XFILLER_126_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15135_ _16509_/Q _15241_/B _15135_/C vssd1 vssd1 vccd1 vccd1 _15135_/X sky130_fd_sc_hd__and3_1
X_12347_ _16099_/Q _12347_/B _12352_/C vssd1 vssd1 vccd1 vccd1 _12347_/Y sky130_fd_sc_hd__nand3_1
XFILLER_142_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15066_ _15066_/A vssd1 vssd1 vccd1 vccd1 _16495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12278_ _13407_/A vssd1 vssd1 vccd1 vccd1 _12501_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_141_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14017_ _16337_/Q _14179_/B _14017_/C vssd1 vssd1 vccd1 vccd1 _14017_/X sky130_fd_sc_hd__and3_1
X_11229_ _16564_/Q vssd1 vssd1 vccd1 vccd1 _11246_/C sky130_fd_sc_hd__inv_2
XFILLER_122_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15968_ _16005_/CLK _15968_/D vssd1 vssd1 vccd1 vccd1 _15968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14919_ _14917_/Y _14918_/X _14914_/C _14915_/C vssd1 vssd1 vccd1 vccd1 _14921_/B
+ sky130_fd_sc_hd__o211ai_1
X_15899_ _16553_/Q _15899_/D vssd1 vssd1 vccd1 vccd1 _15899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ _08440_/A _08339_/A vssd1 vssd1 vccd1 vccd1 _08441_/B sky130_fd_sc_hd__or2b_1
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08371_ _08371_/A _08244_/A vssd1 vssd1 vccd1 vccd1 _08377_/B sky130_fd_sc_hd__or2b_1
XFILLER_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09825_ _11828_/A vssd1 vssd1 vccd1 vccd1 _10300_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09756_ _09756_/A vssd1 vssd1 vccd1 vccd1 _09756_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08707_ _10430_/A vssd1 vssd1 vccd1 vccd1 _15338_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09687_/A _09687_/B vssd1 vssd1 vccd1 vccd1 _09687_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _14821_/A vssd1 vssd1 vccd1 vccd1 _10755_/B sky130_fd_sc_hd__clkbuf_4
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _08567_/X _08568_/X _08565_/X _15367_/B vssd1 vssd1 vccd1 vccd1 _15453_/D
+ sky130_fd_sc_hd__a31oi_1
XFILLER_23_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10600_ _15845_/Q _10646_/B _10606_/C vssd1 vssd1 vccd1 vccd1 _10600_/Y sky130_fd_sc_hd__nand3_1
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ _15992_/Q _11750_/B _11586_/C vssd1 vssd1 vccd1 vccd1 _11582_/C sky130_fd_sc_hd__nand3_1
XFILLER_23_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10531_ _10536_/C vssd1 vssd1 vccd1 vccd1 _10546_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13250_ _16228_/Q _13305_/B _13250_/C vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__and3_1
XFILLER_10_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10462_ _15821_/Q _10463_/C _10360_/X vssd1 vssd1 vccd1 vccd1 _10464_/A sky130_fd_sc_hd__a21oi_1
XFILLER_108_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ _12222_/A _12201_/B _12201_/C vssd1 vssd1 vccd1 vccd1 _12202_/A sky130_fd_sc_hd__and3_1
XFILLER_108_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _13190_/A _13181_/B _13181_/C vssd1 vssd1 vccd1 vccd1 _13182_/A sky130_fd_sc_hd__and3_1
X_10393_ _10393_/A vssd1 vssd1 vccd1 vccd1 _10393_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12132_ _13545_/A vssd1 vssd1 vccd1 vccd1 _13264_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_124_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12063_ _12084_/A _12063_/B _12067_/B vssd1 vssd1 vccd1 vccd1 _16059_/D sky130_fd_sc_hd__nor3_1
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11014_ _11014_/A _11014_/B _11014_/C vssd1 vssd1 vccd1 vccd1 _11015_/C sky130_fd_sc_hd__nand3_1
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15822_ _16551_/CLK _15822_/D vssd1 vssd1 vccd1 vccd1 _15822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15753_ _15791_/CLK _15753_/D vssd1 vssd1 vccd1 vccd1 _15753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ _13377_/A vssd1 vssd1 vccd1 vccd1 _13080_/A sky130_fd_sc_hd__buf_2
X_14704_ _16438_/Q _14875_/B _14710_/C vssd1 vssd1 vccd1 vccd1 _14704_/Y sky130_fd_sc_hd__nand3_1
X_11916_ _16040_/Q _12031_/B _11922_/C vssd1 vssd1 vccd1 vccd1 _11918_/C sky130_fd_sc_hd__nand3_1
X_15684_ _15791_/CLK _15684_/D vssd1 vssd1 vccd1 vccd1 _15684_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _16177_/Q _13009_/B _12896_/C vssd1 vssd1 vccd1 vccd1 _12896_/Y sky130_fd_sc_hd__nand3_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14635_ _14629_/C _14630_/C _14632_/Y _14633_/X vssd1 vssd1 vccd1 vccd1 _14636_/C
+ sky130_fd_sc_hd__a211o_1
X_11847_ _11901_/A _11852_/C vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__or2_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14566_ _14624_/A _14566_/B _14571_/A vssd1 vssd1 vccd1 vccd1 _16416_/D sky130_fd_sc_hd__nor3_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _16020_/Q _11785_/C _11719_/X vssd1 vssd1 vccd1 vccd1 _11778_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13517_ _13526_/A _13517_/B _13517_/C vssd1 vssd1 vccd1 vccd1 _13518_/A sky130_fd_sc_hd__and3_1
X_16305_ _16346_/CLK _16305_/D vssd1 vssd1 vccd1 vccd1 _16305_/Q sky130_fd_sc_hd__dfxtp_1
X_10729_ _15871_/Q _10729_/B _10735_/C vssd1 vssd1 vccd1 vccd1 _10731_/C sky130_fd_sc_hd__nand3_1
X_14497_ _14535_/A _14497_/B _14497_/C vssd1 vssd1 vccd1 vccd1 _14498_/A sky130_fd_sc_hd__and3_1
XFILLER_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16236_ _16237_/CLK _16236_/D vssd1 vssd1 vccd1 vccd1 _16236_/Q sky130_fd_sc_hd__dfxtp_1
X_13448_ _13470_/A _13448_/B _13448_/C vssd1 vssd1 vccd1 vccd1 _13449_/A sky130_fd_sc_hd__and3_1
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ _16237_/CLK _16167_/D vssd1 vssd1 vccd1 vccd1 _16167_/Q sky130_fd_sc_hd__dfxtp_1
X_13379_ _13393_/C vssd1 vssd1 vccd1 vccd1 _13401_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15118_ _15152_/A _15118_/B _15118_/C vssd1 vssd1 vccd1 vccd1 _15119_/A sky130_fd_sc_hd__and3_1
X_16098_ _16118_/CLK _16098_/D vssd1 vssd1 vccd1 vccd1 _16098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15049_ _16494_/Q _15261_/B _15049_/C vssd1 vssd1 vccd1 vccd1 _15057_/A sky130_fd_sc_hd__and3_1
X_07940_ _08265_/A _07939_/B _07939_/C vssd1 vssd1 vccd1 vccd1 _07941_/B sky130_fd_sc_hd__a21oi_1
XFILLER_141_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07871_ _16478_/Q _16460_/Q vssd1 vssd1 vccd1 vccd1 _07872_/B sky130_fd_sc_hd__nand2_1
XFILLER_122_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09610_ _09655_/A _09610_/B vssd1 vssd1 vccd1 vccd1 _09611_/B sky130_fd_sc_hd__and2_1
XFILLER_83_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09541_ _15646_/Q _09669_/B _09541_/C vssd1 vssd1 vccd1 vccd1 _09546_/A sky130_fd_sc_hd__and3_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09472_ _15632_/Q _09472_/B _09472_/C vssd1 vssd1 vccd1 vccd1 _09472_/X sky130_fd_sc_hd__and3_1
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ _08419_/X _08421_/X _08422_/Y vssd1 vssd1 vccd1 vccd1 _15448_/D sky130_fd_sc_hd__o21a_1
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ _08354_/A _08354_/B vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08285_ _08096_/A _08096_/B _08284_/Y vssd1 vssd1 vccd1 vccd1 _08404_/B sky130_fd_sc_hd__o21a_1
XFILLER_149_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09808_ _09809_/B _09809_/C _09809_/A vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__a21o_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09739_ _15686_/Q _09966_/B _09739_/C vssd1 vssd1 vccd1 vccd1 _09739_/X sky130_fd_sc_hd__and3_1
XFILLER_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _12748_/A _12748_/B _12749_/X vssd1 vssd1 vccd1 vccd1 _16156_/D sky130_fd_sc_hd__a21oi_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11717_/A _11701_/B _11701_/C vssd1 vssd1 vccd1 vccd1 _11702_/A sky130_fd_sc_hd__and3_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12681_/A _12681_/B _12681_/C vssd1 vssd1 vccd1 vccd1 _12682_/A sky130_fd_sc_hd__and3_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _16395_/Q _14472_/B _14427_/C vssd1 vssd1 vccd1 vccd1 _14420_/X sky130_fd_sc_hd__and3_1
X_11632_ _16000_/Q _11750_/B _11638_/C vssd1 vssd1 vccd1 vccd1 _11634_/C sky130_fd_sc_hd__nand3_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14351_ _16385_/Q _14458_/B _14351_/C vssd1 vssd1 vccd1 vccd1 _14351_/X sky130_fd_sc_hd__and3_1
XFILLER_7_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11563_ _11563_/A _11563_/B vssd1 vssd1 vccd1 vccd1 _11569_/C sky130_fd_sc_hd__nor2_1
XFILLER_11_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _13302_/A _13302_/B _13302_/C vssd1 vssd1 vccd1 vccd1 _13303_/A sky130_fd_sc_hd__and3_1
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ _10563_/A _10514_/B _10519_/B vssd1 vssd1 vccd1 vccd1 _15827_/D sky130_fd_sc_hd__nor3_1
X_14282_ _14317_/C vssd1 vssd1 vccd1 vccd1 _14323_/C sky130_fd_sc_hd__clkbuf_2
X_11494_ _15980_/Q _11607_/B _11494_/C vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__and3_1
X_16021_ _16554_/Q _16021_/D vssd1 vssd1 vccd1 vccd1 _16021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13233_ _16226_/Q _13235_/C _13006_/X vssd1 vssd1 vccd1 vccd1 _13233_/Y sky130_fd_sc_hd__a21oi_1
X_10445_ _15819_/Q _10457_/C _10393_/X vssd1 vssd1 vccd1 vccd1 _10445_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ _16216_/Q _13164_/B _13171_/C vssd1 vssd1 vccd1 vccd1 _13166_/C sky130_fd_sc_hd__nand3_1
X_10376_ _10388_/C vssd1 vssd1 vccd1 vccd1 _10402_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12115_ _14220_/A vssd1 vssd1 vccd1 vccd1 _12683_/A sky130_fd_sc_hd__clkbuf_2
X_13095_ _13095_/A vssd1 vssd1 vccd1 vccd1 _16205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12046_ _12043_/Y _12044_/X _12045_/Y _12041_/C vssd1 vssd1 vccd1 vccd1 _12048_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _16595_/CLK _15805_/D vssd1 vssd1 vccd1 vccd1 _15805_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13997_ _13997_/A _13997_/B _13997_/C vssd1 vssd1 vccd1 vccd1 _13998_/C sky130_fd_sc_hd__or3_1
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15736_ _15812_/CLK _15736_/D vssd1 vssd1 vccd1 vccd1 _15736_/Q sky130_fd_sc_hd__dfxtp_1
X_12948_ _12963_/A _12948_/B _12948_/C vssd1 vssd1 vccd1 vccd1 _12949_/A sky130_fd_sc_hd__and3_1
XFILLER_61_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15667_ _15791_/CLK _15667_/D vssd1 vssd1 vccd1 vccd1 _15667_/Q sky130_fd_sc_hd__dfxtp_1
X_12879_ _13443_/A vssd1 vssd1 vccd1 vccd1 _12879_/X sky130_fd_sc_hd__buf_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14618_ _14633_/C vssd1 vssd1 vccd1 vccd1 _14640_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15598_ _16551_/CLK _15598_/D vssd1 vssd1 vccd1 vccd1 _15598_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14549_ _14549_/A _14549_/B vssd1 vssd1 vccd1 vccd1 _14550_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08070_ _16487_/Q vssd1 vssd1 vccd1 vccd1 _14902_/A sky130_fd_sc_hd__inv_2
XFILLER_134_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16219_ _16237_/CLK _16219_/D vssd1 vssd1 vccd1 vccd1 _16219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08972_ _15530_/Q _08991_/C _08843_/X vssd1 vssd1 vccd1 vccd1 _08974_/B sky130_fd_sc_hd__a21oi_1
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16677__82 vssd1 vssd1 vccd1 vccd1 _16677__82/HI _16753_/A sky130_fd_sc_hd__conb_1
X_07923_ _13603_/A _07923_/B vssd1 vssd1 vccd1 vccd1 _07932_/A sky130_fd_sc_hd__xnor2_1
XFILLER_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07854_ _15480_/Q vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__inv_2
X_07785_ _07787_/A vssd1 vssd1 vccd1 vccd1 _07785_/Y sky130_fd_sc_hd__inv_2
X_09524_ _09744_/A vssd1 vssd1 vccd1 vccd1 _09524_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09455_ _09455_/A vssd1 vssd1 vccd1 vccd1 _15626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08406_ _08473_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08407_/B sky130_fd_sc_hd__xor2_1
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09386_ _09381_/Y _09385_/X _09304_/X vssd1 vssd1 vccd1 vccd1 _09386_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08337_ _08443_/A _08337_/B vssd1 vssd1 vccd1 vccd1 _08338_/B sky130_fd_sc_hd__nand2_2
XFILLER_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08268_ _08268_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08386_/B sky130_fd_sc_hd__xnor2_1
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08199_ _08020_/A _08197_/Y _08198_/Y vssd1 vssd1 vccd1 vccd1 _08227_/A sky130_fd_sc_hd__a21o_2
X_10230_ _10235_/C vssd1 vssd1 vccd1 vccd1 _10247_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10161_ _10161_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10162_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10092_ _15756_/Q _10300_/C _10099_/C vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__and3_1
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13920_ _16324_/Q _13929_/C _13698_/X vssd1 vssd1 vccd1 vccd1 _13920_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13851_ _13866_/A _13851_/B _13851_/C vssd1 vssd1 vccd1 vccd1 _13852_/A sky130_fd_sc_hd__and3_1
XFILLER_28_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12802_ _12802_/A _12802_/B vssd1 vssd1 vccd1 vccd1 _12808_/C sky130_fd_sc_hd__nor2_1
XFILLER_62_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13782_ _16303_/Q _13822_/C _13781_/X vssd1 vssd1 vccd1 vccd1 _13784_/B sky130_fd_sc_hd__a21oi_1
X_16570_ _16570_/CLK _16570_/D vssd1 vssd1 vccd1 vccd1 _16570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10994_ _10994_/A _10994_/B vssd1 vssd1 vccd1 vccd1 _10995_/B sky130_fd_sc_hd__nor2_1
X_12733_ _16154_/Q _12904_/B _12739_/C vssd1 vssd1 vccd1 vccd1 _12733_/Y sky130_fd_sc_hd__nand3_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15521_ _16551_/CLK _15521_/D vssd1 vssd1 vccd1 vccd1 _15521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _16570_/CLK _15452_/D vssd1 vssd1 vccd1 vccd1 _15452_/Q sky130_fd_sc_hd__dfxtp_1
X_12664_ _12662_/Y _12663_/X _12659_/C _12660_/C vssd1 vssd1 vccd1 vccd1 _12666_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14424_/A _14403_/B _14403_/C vssd1 vssd1 vccd1 vccd1 _14404_/A sky130_fd_sc_hd__and3_1
X_11615_ _11615_/A _11615_/B vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__nor2_1
X_15383_ _15989_/Q _15988_/Q _15987_/Q _15378_/X vssd1 vssd1 vccd1 vccd1 _16569_/D
+ sky130_fd_sc_hd__o31a_1
X_12595_ _13725_/A vssd1 vssd1 vccd1 vccd1 _12818_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ _14334_/A vssd1 vssd1 vccd1 vccd1 _16381_/D sky130_fd_sc_hd__clkbuf_1
X_11546_ _11544_/Y _11539_/C _11541_/Y _11542_/X vssd1 vssd1 vccd1 vccd1 _11547_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14265_ _14828_/A vssd1 vssd1 vccd1 vccd1 _14265_/X sky130_fd_sc_hd__clkbuf_2
X_11477_ _11477_/A vssd1 vssd1 vccd1 vccd1 _15976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16004_ _16005_/CLK _16004_/D vssd1 vssd1 vccd1 vccd1 _16004_/Q sky130_fd_sc_hd__dfxtp_1
X_13216_ _14060_/A vssd1 vssd1 vccd1 vccd1 _13216_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10428_ _15816_/Q _10483_/B _10428_/C vssd1 vssd1 vccd1 vccd1 _10436_/A sky130_fd_sc_hd__and3_1
X_14196_ _14194_/Y _14190_/C _14192_/Y _14193_/X vssd1 vssd1 vccd1 vccd1 _14197_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13315_/A _13151_/C vssd1 vssd1 vccd1 vccd1 _13147_/X sky130_fd_sc_hd__or2_1
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _10429_/A _10359_/B _10364_/B vssd1 vssd1 vccd1 vccd1 _15800_/D sky130_fd_sc_hd__nor3_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13074_/Y _13084_/A _13077_/Y _13072_/C vssd1 vssd1 vccd1 vccd1 _13080_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12029_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12029_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15719_ _15812_/CLK _15719_/D vssd1 vssd1 vccd1 vccd1 _15719_/Q sky130_fd_sc_hd__dfxtp_1
X_16699_ _16699_/A _07798_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_34_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09240_ _09240_/A _09244_/C vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__and2_1
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ _09400_/A vssd1 vssd1 vccd1 vccd1 _09256_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08122_ _10379_/C _07894_/B _08121_/Y vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__o21ai_2
XFILLER_147_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08053_ _11004_/A _08053_/B vssd1 vssd1 vccd1 vccd1 _08094_/A sky130_fd_sc_hd__xnor2_4
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08955_ _08949_/B _08952_/B _08914_/X vssd1 vssd1 vccd1 vccd1 _08963_/C sky130_fd_sc_hd__o21a_1
XFILLER_102_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07906_ _16601_/Q vssd1 vssd1 vccd1 vccd1 _13322_/A sky130_fd_sc_hd__clkinv_2
XFILLER_56_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08886_ _09126_/A vssd1 vssd1 vccd1 vccd1 _09756_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07837_ _07837_/A vssd1 vssd1 vccd1 vccd1 _07842_/A sky130_fd_sc_hd__buf_12
XFILLER_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07768_ _07768_/A vssd1 vssd1 vccd1 vccd1 _07768_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _15639_/Q _09636_/B _09507_/C vssd1 vssd1 vccd1 vccd1 _09513_/A sky130_fd_sc_hd__and3_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _10469_/A vssd1 vssd1 vccd1 vccd1 _09438_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _10294_/C vssd1 vssd1 vccd1 vccd1 _09369_/X sky130_fd_sc_hd__buf_2
XFILLER_40_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11400_ _11436_/C vssd1 vssd1 vccd1 vccd1 _11444_/C sky130_fd_sc_hd__clkbuf_2
X_12380_ _16105_/Q _12487_/B _12380_/C vssd1 vssd1 vccd1 vccd1 _12380_/X sky130_fd_sc_hd__and3_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ _11331_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11336_/C sky130_fd_sc_hd__nor2_1
XFILLER_119_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14050_ _14160_/A vssd1 vssd1 vccd1 vccd1 _14090_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11262_ _11258_/Y _11259_/X _11261_/Y _11256_/C vssd1 vssd1 vccd1 vccd1 _11264_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_106_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13001_ _16193_/Q _13053_/B _13001_/C vssd1 vssd1 vccd1 vccd1 _13001_/X sky130_fd_sc_hd__and3_1
X_10213_ _11150_/A vssd1 vssd1 vccd1 vccd1 _10463_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11193_ _11208_/A _11193_/B _11193_/C vssd1 vssd1 vccd1 vccd1 _11194_/A sky130_fd_sc_hd__and3_1
XFILLER_134_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10144_ _10142_/Y _10136_/C _10139_/Y _10140_/X vssd1 vssd1 vccd1 vccd1 _10145_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10075_ _15753_/Q _10106_/C _09943_/X vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__a21oi_1
X_14952_ _14950_/A _14950_/B _14951_/X vssd1 vssd1 vccd1 vccd1 _16476_/D sky130_fd_sc_hd__a21oi_1
XFILLER_48_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13903_ _13918_/A _13903_/B _13903_/C vssd1 vssd1 vccd1 vccd1 _13904_/A sky130_fd_sc_hd__and3_1
X_14883_ _14880_/Y _14889_/A _14882_/Y _14878_/C vssd1 vssd1 vccd1 vccd1 _14885_/B
+ sky130_fd_sc_hd__o211a_1
X_13834_ _16610_/Q vssd1 vssd1 vccd1 vccd1 _13848_/C sky130_fd_sc_hd__clkinv_2
XFILLER_16_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16553_ _16554_/Q _16553_/D vssd1 vssd1 vccd1 vccd1 _16553_/Q sky130_fd_sc_hd__dfxtp_4
X_13765_ _16301_/Q _13929_/B _13765_/C vssd1 vssd1 vccd1 vccd1 _13774_/B sky130_fd_sc_hd__and3_1
X_10977_ _11828_/A vssd1 vssd1 vccd1 vccd1 _11205_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _16551_/CLK _15504_/D vssd1 vssd1 vccd1 vccd1 _15504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12716_ _12716_/A vssd1 vssd1 vccd1 vccd1 _16151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16484_ _16607_/CLK _16484_/D vssd1 vssd1 vccd1 vccd1 _16484_/Q sky130_fd_sc_hd__dfxtp_1
X_13696_ _13696_/A _13696_/B _13696_/C vssd1 vssd1 vccd1 vccd1 _13697_/A sky130_fd_sc_hd__and3_1
X_12647_ _12663_/C vssd1 vssd1 vccd1 vccd1 _12670_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15435_ _16317_/Q _16316_/Q _16315_/Q _15434_/X vssd1 vssd1 vccd1 vccd1 _16610_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15366_ _16554_/Q _15366_/B vssd1 vssd1 vccd1 vccd1 _16554_/D sky130_fd_sc_hd__nor2_1
X_12578_ _16133_/Q _12798_/B _12578_/C vssd1 vssd1 vccd1 vccd1 _12586_/B sky130_fd_sc_hd__and3_1
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11529_ _15985_/Q _11638_/B _11529_/C vssd1 vssd1 vccd1 vccd1 _11529_/X sky130_fd_sc_hd__and3_1
X_14317_ _16380_/Q _14427_/B _14317_/C vssd1 vssd1 vccd1 vccd1 _14325_/A sky130_fd_sc_hd__and3_1
X_15297_ _16708_/A _15306_/A vssd1 vssd1 vccd1 vccd1 _15299_/B sky130_fd_sc_hd__and2_1
XFILLER_144_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14248_ _14256_/A _14248_/B _14248_/C vssd1 vssd1 vccd1 vccd1 _14249_/A sky130_fd_sc_hd__and3_1
XFILLER_132_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14179_ _16361_/Q _14179_/B _14179_/C vssd1 vssd1 vccd1 vccd1 _14179_/X sky130_fd_sc_hd__and3_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16647__52 vssd1 vssd1 vccd1 vccd1 _16647__52/HI _16723_/A sky130_fd_sc_hd__conb_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08740_ _08733_/B _08736_/B _08698_/X vssd1 vssd1 vccd1 vccd1 _08752_/C sky130_fd_sc_hd__o21a_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08671_ input9/X vssd1 vssd1 vccd1 vccd1 _14848_/A sky130_fd_sc_hd__buf_4
XFILLER_54_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ _09367_/A _09223_/B _09223_/C vssd1 vssd1 vccd1 vccd1 _09224_/A sky130_fd_sc_hd__and3_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09154_ _09849_/A _09154_/B vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__or2_1
XFILLER_148_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08105_ _08110_/A _08111_/B vssd1 vssd1 vccd1 vccd1 _08106_/B sky130_fd_sc_hd__xnor2_2
XFILLER_108_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09085_ _08923_/X _09083_/A _09039_/X vssd1 vssd1 vccd1 vccd1 _09086_/B sky130_fd_sc_hd__o21ai_1
XFILLER_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08036_ _14444_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _08038_/B sky130_fd_sc_hd__xnor2_1
XFILLER_150_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09987_ _15736_/Q _10285_/C _09987_/C vssd1 vssd1 vccd1 vccd1 _09994_/A sky130_fd_sc_hd__and3_1
XFILLER_89_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08938_ _08939_/B _08939_/C _08939_/A vssd1 vssd1 vccd1 vccd1 _08940_/B sky130_fd_sc_hd__a21o_1
XFILLER_123_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08869_ _08869_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08870_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10900_ _15896_/Q _10900_/B _10907_/C vssd1 vssd1 vccd1 vccd1 _10902_/C sky130_fd_sc_hd__nand3_1
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11880_ _11878_/Y _11872_/C _11876_/Y _11877_/X vssd1 vssd1 vccd1 vccd1 _11881_/C
+ sky130_fd_sc_hd__a211o_1
X_10831_ _10868_/C vssd1 vssd1 vccd1 vccd1 _10878_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ _13550_/A vssd1 vssd1 vccd1 vccd1 _16269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10762_ _15353_/A _10762_/B vssd1 vssd1 vccd1 vccd1 _10762_/Y sky130_fd_sc_hd__nor2_1
Xrepeater16 _16555_/Q vssd1 vssd1 vccd1 vccd1 _16261_/CLK sky130_fd_sc_hd__buf_12
XFILLER_16_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12501_ _16123_/Q _12501_/B _12510_/C vssd1 vssd1 vccd1 vccd1 _12501_/X sky130_fd_sc_hd__and3_1
X_13481_ _13481_/A _13481_/B vssd1 vssd1 vccd1 vccd1 _13482_/B sky130_fd_sc_hd__nor2_1
X_10693_ _10690_/Y _10691_/X _10692_/Y _10688_/C vssd1 vssd1 vccd1 vccd1 _10695_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15220_ _15218_/A _15218_/B _15219_/X vssd1 vssd1 vccd1 vccd1 _16521_/D sky130_fd_sc_hd__a21oi_1
X_12432_ _12453_/A _12432_/B _12432_/C vssd1 vssd1 vccd1 vccd1 _12433_/A sky130_fd_sc_hd__and3_1
XFILLER_139_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15151_ _15149_/Y _15145_/C _15147_/Y _15148_/X vssd1 vssd1 vccd1 vccd1 _15152_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _12363_/A vssd1 vssd1 vccd1 vccd1 _16101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _14102_/A _14110_/B vssd1 vssd1 vccd1 vccd1 _14104_/A sky130_fd_sc_hd__or2_1
X_11314_ _15955_/Q _11322_/C _11202_/X vssd1 vssd1 vccd1 vccd1 _11314_/Y sky130_fd_sc_hd__a21oi_1
X_15082_ _16500_/Q _15090_/C _14858_/X vssd1 vssd1 vccd1 vccd1 _15082_/Y sky130_fd_sc_hd__a21oi_1
X_12294_ input6/X vssd1 vssd1 vccd1 vccd1 _13423_/A sky130_fd_sc_hd__buf_2
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14033_ _14030_/Y _14031_/X _14032_/Y _14027_/C vssd1 vssd1 vccd1 vccd1 _14035_/B
+ sky130_fd_sc_hd__o211ai_1
X_11245_ _15945_/Q _11253_/C _11188_/X vssd1 vssd1 vccd1 vccd1 _11245_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _15935_/Q _11217_/C _10951_/X vssd1 vssd1 vccd1 vccd1 _11180_/B sky130_fd_sc_hd__a21oi_1
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10127_ _15763_/Q _10288_/C _10133_/C vssd1 vssd1 vccd1 vccd1 _10129_/C sky130_fd_sc_hd__nand3_1
XFILLER_121_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15984_ _16005_/CLK _15984_/D vssd1 vssd1 vccd1 vccd1 _15984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10058_ _10058_/A _10058_/B vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__or2_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14935_ _14933_/Y _14928_/C _14930_/Y _14931_/X vssd1 vssd1 vccd1 vccd1 _14936_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14866_ _16465_/Q _15033_/B _14867_/C vssd1 vssd1 vccd1 vccd1 _14866_/X sky130_fd_sc_hd__and3_1
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16605_ _16607_/CLK _16605_/D vssd1 vssd1 vccd1 vccd1 _16605_/Q sky130_fd_sc_hd__dfxtp_1
X_13817_ _16307_/Q _14039_/B _13822_/C vssd1 vssd1 vccd1 vccd1 _13817_/Y sky130_fd_sc_hd__nand3_1
XFILLER_91_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14797_ _14797_/A vssd1 vssd1 vccd1 vccd1 _16453_/D sky130_fd_sc_hd__clkbuf_1
X_16536_ _16570_/CLK _16536_/D vssd1 vssd1 vccd1 vccd1 _16705_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13748_ _13756_/A _13748_/B _13748_/C vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__and3_1
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16467_ _16607_/CLK _16467_/D vssd1 vssd1 vccd1 vccd1 _16467_/Q sky130_fd_sc_hd__dfxtp_1
X_13679_ _13696_/A _13679_/B _13679_/C vssd1 vssd1 vccd1 vccd1 _13680_/A sky130_fd_sc_hd__and3_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15418_ _16205_/Q _16204_/Q _16203_/Q _15416_/X vssd1 vssd1 vccd1 vccd1 _16596_/D
+ sky130_fd_sc_hd__o31a_1
X_16398_ input11/X _16398_/D vssd1 vssd1 vccd1 vccd1 _16398_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15349_ _15349_/A _15349_/B vssd1 vssd1 vccd1 vccd1 _15350_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09910_ _09910_/A _09910_/B _09910_/C vssd1 vssd1 vccd1 vccd1 _09911_/C sky130_fd_sc_hd__nand3_1
XFILLER_104_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09841_ _09841_/A _09841_/B _09847_/B vssd1 vssd1 vccd1 vccd1 _15701_/D sky130_fd_sc_hd__nor3_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09772_ _09766_/C _09767_/C _09769_/Y _09776_/A vssd1 vssd1 vccd1 vccd1 _09776_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08723_/A _08723_/B _08723_/C vssd1 vssd1 vccd1 vccd1 _08724_/C sky130_fd_sc_hd__nand3_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08654_ _09615_/A vssd1 vssd1 vccd1 vccd1 _08654_/X sky130_fd_sc_hd__buf_2
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08585_ _15459_/Q _08590_/C _15335_/B vssd1 vssd1 vccd1 vccd1 _08592_/B sky130_fd_sc_hd__a21o_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09206_ _09206_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _15577_/D sky130_fd_sc_hd__nor2_1
XFILLER_10_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09137_ _09148_/A _09137_/B _09141_/A vssd1 vssd1 vccd1 vccd1 _15562_/D sky130_fd_sc_hd__nor3_1
XFILLER_135_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09068_ _09148_/A _09068_/B _09072_/B vssd1 vssd1 vccd1 vccd1 _15546_/D sky130_fd_sc_hd__nor3_1
XFILLER_136_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08019_ _10889_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08197_/A sky130_fd_sc_hd__xnor2_4
XFILLER_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11030_ _11030_/A vssd1 vssd1 vccd1 vccd1 _15913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12981_ _13034_/A vssd1 vssd1 vccd1 vccd1 _13019_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14720_ _14720_/A _14724_/C vssd1 vssd1 vccd1 vccd1 _14720_/X sky130_fd_sc_hd__or2_1
XFILLER_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11932_ _11930_/Y _11925_/C _11927_/Y _11928_/X vssd1 vssd1 vccd1 vccd1 _11933_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11863_ _16032_/Q _12031_/B _11869_/C vssd1 vssd1 vccd1 vccd1 _11865_/C sky130_fd_sc_hd__nand3_1
X_14651_ _14651_/A _14651_/B _14651_/C vssd1 vssd1 vccd1 vccd1 _14652_/A sky130_fd_sc_hd__and3_1
XFILLER_60_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10814_ _10814_/A _10814_/B vssd1 vssd1 vccd1 vccd1 _10816_/B sky130_fd_sc_hd__nor2_1
X_13602_ _13602_/A vssd1 vssd1 vccd1 vccd1 _16277_/D sky130_fd_sc_hd__clkbuf_1
X_14582_ _16420_/Q _14748_/B _14583_/C vssd1 vssd1 vccd1 vccd1 _14582_/X sky130_fd_sc_hd__and3_1
X_11794_ _12924_/A vssd1 vssd1 vccd1 vccd1 _12018_/A sky130_fd_sc_hd__clkbuf_2
X_16321_ _16346_/CLK _16321_/D vssd1 vssd1 vccd1 vccd1 _16321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10745_ _10743_/Y _10738_/C _10741_/Y _10742_/X vssd1 vssd1 vccd1 vccd1 _10746_/C
+ sky130_fd_sc_hd__a211o_1
X_13533_ _16267_/Q _13760_/B _13538_/C vssd1 vssd1 vccd1 vccd1 _13533_/Y sky130_fd_sc_hd__nand3_1
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16252_ _16261_/CLK _16252_/D vssd1 vssd1 vccd1 vccd1 _16252_/Q sky130_fd_sc_hd__dfxtp_1
X_13464_ _14308_/A vssd1 vssd1 vccd1 vccd1 _13464_/X sky130_fd_sc_hd__clkbuf_2
X_10676_ _10676_/A _10676_/B _10681_/A vssd1 vssd1 vccd1 vccd1 _15859_/D sky130_fd_sc_hd__nor3_1
X_15203_ _15200_/Y _15201_/X _15202_/Y _15198_/C vssd1 vssd1 vccd1 vccd1 _15205_/B
+ sky130_fd_sc_hd__o211ai_1
X_12415_ _12468_/A vssd1 vssd1 vccd1 vccd1 _12453_/A sky130_fd_sc_hd__clkbuf_2
X_13395_ _13388_/C _13389_/C _13391_/Y _13393_/X vssd1 vssd1 vccd1 vccd1 _13396_/C
+ sky130_fd_sc_hd__a211o_1
X_16183_ _16237_/CLK _16183_/D vssd1 vssd1 vccd1 vccd1 _16183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15134_ _16509_/Q _15142_/C _10782_/B vssd1 vssd1 vccd1 vccd1 _15134_/Y sky130_fd_sc_hd__a21oi_1
X_12346_ _16100_/Q _12456_/B _12346_/C vssd1 vssd1 vccd1 vccd1 _12354_/A sky130_fd_sc_hd__and3_1
XFILLER_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15065_ _15100_/A _15065_/B _15065_/C vssd1 vssd1 vccd1 vccd1 _15066_/A sky130_fd_sc_hd__and3_1
XFILLER_114_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12277_ input4/X vssd1 vssd1 vccd1 vccd1 _13407_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ _16337_/Q _14024_/C _14015_/X vssd1 vssd1 vccd1 vccd1 _14016_/Y sky130_fd_sc_hd__a21oi_1
X_11228_ _11228_/A vssd1 vssd1 vccd1 vccd1 _15941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11159_ _15933_/Q _11161_/C _11158_/X vssd1 vssd1 vccd1 vccd1 _11162_/A sky130_fd_sc_hd__a21oi_1
XFILLER_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15967_ _16005_/CLK _15967_/D vssd1 vssd1 vccd1 vccd1 _15967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14918_ _16473_/Q _15027_/B _14918_/C vssd1 vssd1 vccd1 vccd1 _14918_/X sky130_fd_sc_hd__and3_1
X_15898_ _16553_/Q _15898_/D vssd1 vssd1 vccd1 vccd1 _15898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14849_ _16462_/Q _15074_/B _14860_/C vssd1 vssd1 vccd1 vccd1 _14855_/A sky130_fd_sc_hd__and3_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _08370_/A _08243_/A vssd1 vssd1 vccd1 vccd1 _08377_/A sky130_fd_sc_hd__or2b_1
X_16519_ _16607_/CLK _16519_/D vssd1 vssd1 vccd1 vccd1 _16519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09824_ _14979_/A vssd1 vssd1 vccd1 vccd1 _11828_/A sky130_fd_sc_hd__buf_8
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09755_ _09755_/A _09755_/B vssd1 vssd1 vccd1 vccd1 _15686_/D sky130_fd_sc_hd__nor2_1
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08706_ _09615_/A vssd1 vssd1 vccd1 vccd1 _08706_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09686_ _15676_/Q _09919_/B _09692_/C vssd1 vssd1 vccd1 vccd1 _09688_/B sky130_fd_sc_hd__and3_1
XFILLER_104_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08637_ _12849_/A vssd1 vssd1 vccd1 vccd1 _14821_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08568_ _15327_/A _08568_/B vssd1 vssd1 vccd1 vccd1 _08568_/X sky130_fd_sc_hd__or2_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ _08538_/A _08499_/B vssd1 vssd1 vccd1 vccd1 _08499_/Y sky130_fd_sc_hd__xnor2_1
X_10530_ _15849_/Q vssd1 vssd1 vccd1 vccd1 _10536_/C sky130_fd_sc_hd__inv_2
XFILLER_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _10563_/A _10461_/B _10465_/B vssd1 vssd1 vccd1 vccd1 _15818_/D sky130_fd_sc_hd__nor3_1
XFILLER_129_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12200_ _12200_/A _12200_/B _12200_/C vssd1 vssd1 vccd1 vccd1 _12201_/C sky130_fd_sc_hd__nand3_1
XFILLER_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13180_ _13178_/Y _13174_/C _13176_/Y _13177_/X vssd1 vssd1 vccd1 vccd1 _13181_/C
+ sky130_fd_sc_hd__a211o_1
X_10392_ _10392_/A vssd1 vssd1 vccd1 vccd1 _15807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12131_ _12185_/A vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12062_ _12060_/Y _12056_/C _12058_/Y _12067_/A vssd1 vssd1 vccd1 vccd1 _12067_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_145_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11013_ _11014_/B _11014_/C _11014_/A vssd1 vssd1 vccd1 vccd1 _11015_/B sky130_fd_sc_hd__a21o_1
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15821_ _16551_/CLK _15821_/D vssd1 vssd1 vccd1 vccd1 _15821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15752_ _15791_/CLK _15752_/D vssd1 vssd1 vccd1 vccd1 _15752_/Q sky130_fd_sc_hd__dfxtp_2
X_12964_ _12964_/A vssd1 vssd1 vccd1 vccd1 _16186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14703_ _16439_/Q _14756_/B _14710_/C vssd1 vssd1 vccd1 vccd1 _14703_/X sky130_fd_sc_hd__and3_1
X_11915_ _16040_/Q _11922_/C _11748_/X vssd1 vssd1 vccd1 vccd1 _11918_/B sky130_fd_sc_hd__a21o_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15791_/CLK _15683_/D vssd1 vssd1 vccd1 vccd1 _15683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _16178_/Q _13059_/B _12896_/C vssd1 vssd1 vccd1 vccd1 _12895_/X sky130_fd_sc_hd__and3_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14634_ _14632_/Y _14633_/X _14629_/C _14630_/C vssd1 vssd1 vccd1 vccd1 _14636_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11846_ _11846_/A _11846_/B vssd1 vssd1 vccd1 vccd1 _11852_/C sky130_fd_sc_hd__nor2_1
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _11777_/A vssd1 vssd1 vccd1 vccd1 _16018_/D sky130_fd_sc_hd__clkbuf_1
X_14565_ _16417_/Q _14790_/B _14576_/C vssd1 vssd1 vccd1 vccd1 _14571_/A sky130_fd_sc_hd__and3_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _16346_/CLK _16304_/D vssd1 vssd1 vccd1 vccd1 _16304_/Q sky130_fd_sc_hd__dfxtp_1
X_10728_ _15871_/Q _10735_/C _09629_/A vssd1 vssd1 vccd1 vccd1 _10731_/B sky130_fd_sc_hd__a21o_1
X_13516_ _13514_/Y _13510_/C _13512_/Y _13513_/X vssd1 vssd1 vccd1 vccd1 _13517_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14496_ _14555_/A _14496_/B _14496_/C vssd1 vssd1 vccd1 vccd1 _14497_/C sky130_fd_sc_hd__or3_1
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16235_ _16237_/CLK _16235_/D vssd1 vssd1 vccd1 vccd1 _16235_/Q sky130_fd_sc_hd__dfxtp_1
X_13447_ _13447_/A _13447_/B _13447_/C vssd1 vssd1 vccd1 vccd1 _13448_/C sky130_fd_sc_hd__nand3_1
X_10659_ _10659_/A _10659_/B vssd1 vssd1 vccd1 vccd1 _10661_/A sky130_fd_sc_hd__or2_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16166_ _16237_/CLK _16166_/D vssd1 vssd1 vccd1 vccd1 _16166_/Q sky130_fd_sc_hd__dfxtp_2
X_13378_ _16602_/Q vssd1 vssd1 vccd1 vccd1 _13393_/C sky130_fd_sc_hd__inv_2
X_15117_ _15117_/A _15117_/B _15117_/C vssd1 vssd1 vccd1 vccd1 _15118_/C sky130_fd_sc_hd__or3_1
XFILLER_126_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12329_ _12329_/A vssd1 vssd1 vccd1 vccd1 _16096_/D sky130_fd_sc_hd__clkbuf_1
X_16097_ _16118_/CLK _16097_/D vssd1 vssd1 vccd1 vccd1 _16097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15048_ _15048_/A vssd1 vssd1 vccd1 vccd1 _15261_/B sky130_fd_sc_hd__buf_2
XFILLER_123_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07870_ _16478_/Q _16460_/Q vssd1 vssd1 vccd1 vccd1 _07872_/A sky130_fd_sc_hd__or2_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09540_ _15646_/Q _09561_/C _09493_/X vssd1 vssd1 vccd1 vccd1 _09542_/B sky130_fd_sc_hd__a21oi_1
XFILLER_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09471_ _09468_/A _09467_/Y _09468_/B vssd1 vssd1 vccd1 vccd1 _09471_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_37_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08422_ _08419_/X _08421_/X _15344_/A vssd1 vssd1 vccd1 vccd1 _08422_/Y sky130_fd_sc_hd__a21oi_1
X_08353_ _08353_/A _08353_/B vssd1 vssd1 vccd1 vccd1 _08365_/A sky130_fd_sc_hd__xor2_4
X_08284_ _15696_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08284_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09807_ _15700_/Q _10288_/C _09816_/C vssd1 vssd1 vccd1 vccd1 _09809_/C sky130_fd_sc_hd__nand3_1
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07999_ _14113_/A _07999_/B vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__xnor2_1
XFILLER_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09738_ _15262_/B vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__buf_2
XFILLER_27_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09669_ _15673_/Q _09669_/B _09669_/C vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__and3_1
XFILLER_55_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11693_/C _11694_/C _11696_/Y _11698_/X vssd1 vssd1 vccd1 vccd1 _11701_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12678_/Y _12673_/C _12675_/Y _12676_/X vssd1 vssd1 vccd1 vccd1 _12681_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _16000_/Q _11638_/C _11463_/X vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__a21o_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _11562_/A _11562_/B vssd1 vssd1 vccd1 vccd1 _11563_/B sky130_fd_sc_hd__nor2_1
X_14350_ _16385_/Q _14358_/C _14294_/X vssd1 vssd1 vccd1 vccd1 _14350_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10513_ _10511_/Y _10506_/C _10508_/Y _10519_/A vssd1 vssd1 vccd1 vccd1 _10519_/B
+ sky130_fd_sc_hd__a211oi_1
X_13301_ _13299_/Y _13295_/C _13297_/Y _13298_/X vssd1 vssd1 vccd1 vccd1 _13302_/C
+ sky130_fd_sc_hd__a211o_1
X_14281_ _14303_/C vssd1 vssd1 vccd1 vccd1 _14317_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11493_ _15980_/Q _11500_/C _11434_/X vssd1 vssd1 vccd1 vccd1 _11493_/Y sky130_fd_sc_hd__a21oi_1
X_13232_ _13232_/A vssd1 vssd1 vccd1 vccd1 _16224_/D sky130_fd_sc_hd__clkbuf_1
X_16020_ _16554_/Q _16020_/D vssd1 vssd1 vccd1 vccd1 _16020_/Q sky130_fd_sc_hd__dfxtp_1
X_10444_ _10444_/A vssd1 vssd1 vccd1 vccd1 _15816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13163_ _16216_/Q _13171_/C _13162_/X vssd1 vssd1 vccd1 vccd1 _13166_/B sky130_fd_sc_hd__a21o_1
X_10375_ _10379_/C vssd1 vssd1 vccd1 vccd1 _10388_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ _12114_/A vssd1 vssd1 vccd1 vccd1 _16066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13094_ _13131_/A _13094_/B _13094_/C vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__and3_1
XFILLER_111_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12045_ _16057_/Q _12160_/B _12045_/C vssd1 vssd1 vccd1 vccd1 _12045_/Y sky130_fd_sc_hd__nand3_1
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15804_ _15812_/CLK _15804_/D vssd1 vssd1 vccd1 vccd1 _15804_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13996_ _13997_/B _13997_/C _13829_/X vssd1 vssd1 vccd1 vccd1 _13998_/B sky130_fd_sc_hd__o21ai_1
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15735_ _16551_/CLK _15735_/D vssd1 vssd1 vccd1 vccd1 _15735_/Q sky130_fd_sc_hd__dfxtp_2
X_12947_ _12941_/C _12942_/C _12944_/Y _12945_/X vssd1 vssd1 vccd1 vccd1 _12948_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_65_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15666_ _15791_/CLK _15666_/D vssd1 vssd1 vccd1 vccd1 _15666_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12936_/A _12878_/B _12883_/A vssd1 vssd1 vccd1 vccd1 _16174_/D sky130_fd_sc_hd__nor3_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14617_ _16442_/Q vssd1 vssd1 vccd1 vccd1 _14633_/C sky130_fd_sc_hd__inv_2
X_11829_ _16026_/Q _12053_/B _11836_/C vssd1 vssd1 vccd1 vccd1 _11829_/Y sky130_fd_sc_hd__nand3_1
X_15597_ _16551_/CLK _15597_/D vssd1 vssd1 vccd1 vccd1 _15597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14548_ _14548_/A _14555_/B vssd1 vssd1 vccd1 vccd1 _14550_/A sky130_fd_sc_hd__or2_1
XFILLER_146_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14479_ _15048_/A vssd1 vssd1 vccd1 vccd1 _14710_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_146_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16218_ _16237_/CLK _16218_/D vssd1 vssd1 vccd1 vccd1 _16218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16149_ _16555_/Q _16149_/D vssd1 vssd1 vccd1 vccd1 _16149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08971_ _08978_/C vssd1 vssd1 vccd1 vccd1 _08991_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_07922_ _07922_/A _07922_/B vssd1 vssd1 vccd1 vccd1 _07923_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07853_ _15447_/Q vssd1 vssd1 vccd1 vccd1 _08108_/A sky130_fd_sc_hd__inv_2
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07784_ _07787_/A vssd1 vssd1 vccd1 vccd1 _07784_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09523_ _09517_/Y _09521_/X _09522_/Y vssd1 vssd1 vccd1 vccd1 _15638_/D sky130_fd_sc_hd__o21a_1
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09454_ _09588_/A _09454_/B _09454_/C vssd1 vssd1 vccd1 vccd1 _09455_/A sky130_fd_sc_hd__and3_1
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08405_ _08287_/A _08287_/B _08404_/Y vssd1 vssd1 vccd1 vccd1 _08473_/B sky130_fd_sc_hd__a21oi_1
X_09385_ _09382_/X _09385_/B vssd1 vssd1 vccd1 vccd1 _09385_/X sky130_fd_sc_hd__and2b_1
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08336_ _08336_/A _08336_/B _08336_/C vssd1 vssd1 vccd1 vccd1 _08337_/B sky130_fd_sc_hd__nand3_1
X_08267_ _08088_/A _08088_/B _08266_/X vssd1 vssd1 vccd1 vccd1 _08268_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08198_ _10889_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08198_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10160_ _10160_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10091_ _15756_/Q _10099_/C _10003_/B vssd1 vssd1 vccd1 vccd1 _10091_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_120_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13850_ _13844_/C _13845_/C _13847_/Y _13848_/X vssd1 vssd1 vccd1 vccd1 _13851_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _12801_/A vssd1 vssd1 vccd1 vccd1 _13032_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13781_ _14060_/A vssd1 vssd1 vccd1 vccd1 _13781_/X sky130_fd_sc_hd__buf_2
X_10993_ _10993_/A _11001_/B vssd1 vssd1 vccd1 vccd1 _10995_/A sky130_fd_sc_hd__or2_1
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15520_ _15791_/CLK _15520_/D vssd1 vssd1 vccd1 vccd1 _15520_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _16155_/Q _12784_/B _12739_/C vssd1 vssd1 vccd1 vccd1 _12732_/X sky130_fd_sc_hd__and3_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _16570_/CLK _15451_/D vssd1 vssd1 vccd1 vccd1 _15451_/Q sky130_fd_sc_hd__dfxtp_1
X_12663_ _16145_/Q _12770_/B _12663_/C vssd1 vssd1 vccd1 vccd1 _12663_/X sky130_fd_sc_hd__and3_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _14402_/A _14402_/B _14402_/C vssd1 vssd1 vccd1 vccd1 _14403_/C sky130_fd_sc_hd__nand3_1
XFILLER_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11614_ _11614_/A _11621_/B vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__or2_1
X_15382_ _15979_/Q _15981_/Q _15980_/Q _15378_/X vssd1 vssd1 vccd1 vccd1 _16568_/D
+ sky130_fd_sc_hd__o31a_1
X_12594_ input9/X vssd1 vssd1 vccd1 vccd1 _13725_/A sky130_fd_sc_hd__buf_2
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14333_ _14369_/A _14333_/B _14333_/C vssd1 vssd1 vccd1 vccd1 _14334_/A sky130_fd_sc_hd__and3_1
XFILLER_128_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11545_ _11541_/Y _11542_/X _11544_/Y _11539_/C vssd1 vssd1 vccd1 vccd1 _11547_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_51_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11476_ _11491_/A _11476_/B _11476_/C vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__and3_1
X_14264_ _14342_/A _14264_/B _14270_/B vssd1 vssd1 vccd1 vccd1 _16371_/D sky130_fd_sc_hd__nor3_1
XFILLER_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16003_ _16005_/CLK _16003_/D vssd1 vssd1 vccd1 vccd1 _16003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10427_ _15816_/Q _10463_/C _10426_/X vssd1 vssd1 vccd1 vccd1 _10429_/B sky130_fd_sc_hd__a21oi_1
X_13215_ _13250_/C vssd1 vssd1 vccd1 vccd1 _13257_/C sky130_fd_sc_hd__clkbuf_2
X_14195_ _14192_/Y _14193_/X _14194_/Y _14190_/C vssd1 vssd1 vccd1 vccd1 _14197_/B
+ sky130_fd_sc_hd__o211ai_1
X_10358_ _10356_/Y _10352_/C _10354_/Y _10364_/A vssd1 vssd1 vccd1 vccd1 _10364_/B
+ sky130_fd_sc_hd__a211oi_1
X_13146_ _13146_/A _13146_/B vssd1 vssd1 vccd1 vccd1 _13151_/C sky130_fd_sc_hd__nor2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _16203_/Q _13194_/B _13082_/C vssd1 vssd1 vccd1 vccd1 _13077_/Y sky130_fd_sc_hd__nand3_1
X_10289_ _10290_/B _10290_/C _10290_/A vssd1 vssd1 vccd1 vccd1 _10291_/B sky130_fd_sc_hd__a21o_1
XFILLER_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12028_ _12084_/A _12028_/B _12033_/A vssd1 vssd1 vccd1 vccd1 _16054_/D sky130_fd_sc_hd__nor3_1
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13979_ _13979_/A vssd1 vssd1 vccd1 vccd1 _13979_/X sky130_fd_sc_hd__buf_2
X_15718_ _15812_/CLK _15718_/D vssd1 vssd1 vccd1 vccd1 _15718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16698_ _16698_/A _07797_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15649_ _15791_/CLK _15649_/D vssd1 vssd1 vccd1 vccd1 _15649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09170_ _15560_/Q _15559_/Q _15558_/Q _09090_/X vssd1 vssd1 vccd1 vccd1 _15570_/D
+ sky130_fd_sc_hd__o31a_1
X_08121_ _15840_/Q _08121_/B vssd1 vssd1 vccd1 vccd1 _08121_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ _11113_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _08053_/B sky130_fd_sc_hd__xnor2_4
XFILLER_127_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08954_ _10112_/A vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07905_ _16599_/Q vssd1 vssd1 vccd1 vccd1 _13212_/A sky130_fd_sc_hd__inv_2
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08885_ _08883_/X _08882_/A _08884_/Y vssd1 vssd1 vccd1 vccd1 _15506_/D sky130_fd_sc_hd__o21a_1
X_07836_ _07836_/A vssd1 vssd1 vccd1 vccd1 _07836_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07767_ _07768_/A vssd1 vssd1 vccd1 vccd1 _07767_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09506_ _15639_/Q _09507_/C _09369_/X vssd1 vssd1 vccd1 vccd1 _09506_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _09291_/X _09435_/B _09436_/Y vssd1 vssd1 vccd1 vccd1 _15621_/D sky130_fd_sc_hd__o21a_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09368_/A vssd1 vssd1 vccd1 vccd1 _15608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08319_ _08319_/A _08145_/A vssd1 vssd1 vccd1 vccd1 _08320_/B sky130_fd_sc_hd__or2b_1
X_09299_ _09749_/A vssd1 vssd1 vccd1 vccd1 _09299_/X sky130_fd_sc_hd__clkbuf_2
X_11330_ _11330_/A _11330_/B vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11261_ _15946_/Q _11488_/B _11268_/C vssd1 vssd1 vccd1 vccd1 _11261_/Y sky130_fd_sc_hd__nand3_1
XFILLER_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10212_ _15776_/Q _10214_/C _10104_/X vssd1 vssd1 vccd1 vccd1 _10215_/A sky130_fd_sc_hd__a21oi_1
X_13000_ _16193_/Q _13009_/C _12887_/X vssd1 vssd1 vccd1 vccd1 _13000_/Y sky130_fd_sc_hd__a21oi_1
X_11192_ _11185_/C _11186_/C _11189_/Y _11190_/X vssd1 vssd1 vccd1 vccd1 _11193_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10143_ _10139_/Y _10140_/X _10142_/Y _10136_/C vssd1 vssd1 vccd1 vccd1 _10145_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_88_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10074_ _10099_/C vssd1 vssd1 vccd1 vccd1 _10106_/C sky130_fd_sc_hd__clkbuf_2
X_14951_ _15005_/A _14956_/C vssd1 vssd1 vccd1 vccd1 _14951_/X sky130_fd_sc_hd__or2_1
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13902_ _13896_/C _13897_/C _13899_/Y _13900_/X vssd1 vssd1 vccd1 vccd1 _13903_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14882_ _16466_/Q _14882_/B _14887_/C vssd1 vssd1 vccd1 vccd1 _14882_/Y sky130_fd_sc_hd__nand3_1
XFILLER_35_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13833_ _13833_/A vssd1 vssd1 vccd1 vccd1 _16309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16552_ _16595_/CLK _16552_/D vssd1 vssd1 vccd1 vccd1 _16702_/A sky130_fd_sc_hd__dfxtp_2
X_13764_ _16301_/Q _13765_/C _13705_/X vssd1 vssd1 vccd1 vccd1 _13766_/A sky130_fd_sc_hd__a21oi_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _15907_/Q _11084_/B _10985_/C vssd1 vssd1 vccd1 vccd1 _10976_/X sky130_fd_sc_hd__and3_1
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15503_ _16570_/CLK _15503_/D vssd1 vssd1 vccd1 vccd1 _15503_/Q sky130_fd_sc_hd__dfxtp_1
X_12715_ _12736_/A _12715_/B _12715_/C vssd1 vssd1 vccd1 vccd1 _12716_/A sky130_fd_sc_hd__and3_1
X_16483_ _16607_/CLK _16483_/D vssd1 vssd1 vccd1 vccd1 _16483_/Q sky130_fd_sc_hd__dfxtp_1
X_13695_ _13693_/Y _13687_/C _13689_/Y _13692_/X vssd1 vssd1 vccd1 vccd1 _13696_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15434_ _15440_/A vssd1 vssd1 vccd1 vccd1 _15434_/X sky130_fd_sc_hd__clkbuf_2
X_12646_ _12646_/A vssd1 vssd1 vccd1 vccd1 _12663_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15365_ _15365_/A _15366_/B vssd1 vssd1 vccd1 vccd1 _16553_/D sky130_fd_sc_hd__nor2_1
X_12577_ _13423_/A vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _16380_/Q _14323_/C _14258_/X vssd1 vssd1 vccd1 vccd1 _14316_/Y sky130_fd_sc_hd__a21oi_1
X_11528_ _15985_/Q _11536_/C _11471_/X vssd1 vssd1 vccd1 vccd1 _11528_/Y sky130_fd_sc_hd__a21oi_1
X_15296_ _15292_/X _15294_/X _15295_/Y vssd1 vssd1 vccd1 vccd1 _16537_/D sky130_fd_sc_hd__o21a_1
X_14247_ _14245_/Y _14240_/C _14242_/Y _14244_/X vssd1 vssd1 vccd1 vccd1 _14248_/C
+ sky130_fd_sc_hd__a211o_1
X_11459_ _15975_/Q _11500_/C _11233_/X vssd1 vssd1 vccd1 vccd1 _11462_/B sky130_fd_sc_hd__a21oi_1
XFILLER_109_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ _16361_/Q _14187_/C _14015_/X vssd1 vssd1 vccd1 vccd1 _14178_/Y sky130_fd_sc_hd__a21oi_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13129_ _13125_/Y _13127_/X _13128_/Y _13123_/C vssd1 vssd1 vccd1 vccd1 _13131_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08670_ _15467_/Q _08689_/C _08576_/X vssd1 vssd1 vccd1 vccd1 _08676_/B sky130_fd_sc_hd__a21oi_1
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16662__67 vssd1 vssd1 vccd1 vccd1 _16662__67/HI _16738_/A sky130_fd_sc_hd__conb_1
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09222_ _09222_/A _09222_/B _09222_/C vssd1 vssd1 vccd1 vccd1 _09223_/C sky130_fd_sc_hd__nand3_1
XFILLER_148_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _09153_/A _09153_/B vssd1 vssd1 vccd1 vccd1 _09154_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08104_ _15069_/A _08104_/B vssd1 vssd1 vccd1 vccd1 _08111_/B sky130_fd_sc_hd__xnor2_2
X_09084_ _09124_/A _09124_/B _09084_/C vssd1 vssd1 vccd1 vccd1 _09086_/A sky130_fd_sc_hd__and3_1
X_08035_ _10332_/C _08035_/B vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__xnor2_4
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09986_ _15736_/Q _10009_/C _09943_/X vssd1 vssd1 vccd1 vccd1 _09988_/B sky130_fd_sc_hd__a21oi_1
XFILLER_77_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08937_ _15522_/Q _09016_/B _08937_/C vssd1 vssd1 vccd1 vccd1 _08939_/C sky130_fd_sc_hd__nand3_1
XFILLER_85_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08868_ _08868_/A _08868_/B vssd1 vssd1 vccd1 vccd1 _08869_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07819_ _07837_/A vssd1 vssd1 vccd1 vccd1 _07824_/A sky130_fd_sc_hd__buf_12
XFILLER_123_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08799_ _15479_/Q _15478_/Q _15477_/Q _08667_/X vssd1 vssd1 vccd1 vccd1 _15489_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_38_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10830_ _10852_/C vssd1 vssd1 vccd1 vccd1 _10868_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10761_ _10756_/B _10759_/B _08705_/B vssd1 vssd1 vccd1 vccd1 _10762_/B sky130_fd_sc_hd__o21a_1
Xrepeater17 _16346_/CLK vssd1 vssd1 vccd1 vccd1 _16389_/CLK sky130_fd_sc_hd__buf_12
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _16123_/Q _12510_/C _12337_/X vssd1 vssd1 vccd1 vccd1 _12500_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ _15863_/Q _10743_/B _10701_/C vssd1 vssd1 vccd1 vccd1 _10692_/Y sky130_fd_sc_hd__nand3_1
X_13480_ _13480_/A _13488_/B vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__or2_1
XFILLER_9_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12431_ _12431_/A _12431_/B _12431_/C vssd1 vssd1 vccd1 vccd1 _12432_/C sky130_fd_sc_hd__nand3_1
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15150_ _15147_/Y _15148_/X _15149_/Y _15145_/C vssd1 vssd1 vccd1 vccd1 _15152_/B
+ sky130_fd_sc_hd__o211ai_1
X_12362_ _12398_/A _12362_/B _12362_/C vssd1 vssd1 vccd1 vccd1 _12363_/A sky130_fd_sc_hd__and3_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14101_ _16349_/Q _14207_/B _14101_/C vssd1 vssd1 vccd1 vccd1 _14110_/B sky130_fd_sc_hd__and3_1
XFILLER_138_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11313_ _11313_/A vssd1 vssd1 vccd1 vccd1 _15953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12293_ _16093_/Q _12296_/C _12292_/X vssd1 vssd1 vccd1 vccd1 _12297_/A sky130_fd_sc_hd__a21oi_1
X_15081_ _15081_/A vssd1 vssd1 vccd1 vccd1 _16498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11244_ _11244_/A vssd1 vssd1 vccd1 vccd1 _15943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14032_ _16338_/Q _14032_/B _14038_/C vssd1 vssd1 vccd1 vccd1 _14032_/Y sky130_fd_sc_hd__nand3_1
XFILLER_122_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11175_ _11211_/C vssd1 vssd1 vccd1 vccd1 _11217_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10126_ _15763_/Q _10133_/C _10729_/B vssd1 vssd1 vccd1 vccd1 _10129_/B sky130_fd_sc_hd__a21o_1
X_15983_ _16005_/CLK _15983_/D vssd1 vssd1 vccd1 vccd1 _15983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10057_ _15749_/Q _10313_/C _10057_/C vssd1 vssd1 vccd1 vccd1 _10058_/B sky130_fd_sc_hd__and3_1
X_14934_ _14930_/Y _14931_/X _14933_/Y _14928_/C vssd1 vssd1 vccd1 vccd1 _14936_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_94_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14865_ _16465_/Q _14867_/C _14694_/X vssd1 vssd1 vccd1 vccd1 _14865_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16604_ _16607_/CLK _16604_/D vssd1 vssd1 vccd1 vccd1 _16604_/Q sky130_fd_sc_hd__dfxtp_1
X_13816_ _14095_/A vssd1 vssd1 vccd1 vccd1 _14039_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14796_ _14819_/A _14796_/B _14796_/C vssd1 vssd1 vccd1 vccd1 _14797_/A sky130_fd_sc_hd__and3_1
X_16535_ _16570_/CLK _16535_/D vssd1 vssd1 vccd1 vccd1 _16704_/A sky130_fd_sc_hd__dfxtp_1
X_13747_ _13745_/Y _13741_/C _13743_/Y _13744_/X vssd1 vssd1 vccd1 vccd1 _13748_/C
+ sky130_fd_sc_hd__a211o_1
X_10959_ _10959_/A _10959_/B _10959_/C vssd1 vssd1 vccd1 vccd1 _10960_/C sky130_fd_sc_hd__nand3_1
XFILLER_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16466_ _16607_/CLK _16466_/D vssd1 vssd1 vccd1 vccd1 _16466_/Q sky130_fd_sc_hd__dfxtp_1
X_13678_ _13670_/C _13671_/C _13673_/Y _13676_/X vssd1 vssd1 vccd1 vccd1 _13679_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15417_ _16197_/Q _16196_/Q _16195_/Q _15416_/X vssd1 vssd1 vccd1 vccd1 _16595_/D
+ sky130_fd_sc_hd__o31a_1
X_12629_ _16139_/Q _12629_/B _12634_/C vssd1 vssd1 vccd1 vccd1 _12629_/Y sky130_fd_sc_hd__nand3_1
X_16397_ input11/X _16397_/D vssd1 vssd1 vccd1 vccd1 _16397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15348_ _15348_/A _15348_/B vssd1 vssd1 vccd1 vccd1 _15349_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15279_ _16450_/Q _16449_/Q _16448_/Q _15172_/X vssd1 vssd1 vccd1 vccd1 _16534_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_145_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09840_ _09838_/Y _09831_/C _09835_/Y _09847_/A vssd1 vssd1 vccd1 vccd1 _09847_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ _09769_/Y _09776_/A _09766_/C _09767_/C vssd1 vssd1 vccd1 vccd1 _09773_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _08723_/B _08723_/C _08723_/A vssd1 vssd1 vccd1 vccd1 _08724_/B sky130_fd_sc_hd__a21o_1
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08653_ _09898_/A vssd1 vssd1 vccd1 vccd1 _09615_/A sky130_fd_sc_hd__buf_2
XFILLER_82_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _09056_/A vssd1 vssd1 vccd1 vccd1 _15335_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09205_ _09125_/X _09203_/A _09126_/X vssd1 vssd1 vccd1 vccd1 _09206_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09136_ _15566_/Q _15332_/B _09139_/C vssd1 vssd1 vccd1 vccd1 _09141_/A sky130_fd_sc_hd__and3_1
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09067_ _09059_/C _09060_/C _09064_/Y _09072_/A vssd1 vssd1 vccd1 vccd1 _09072_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08018_ _12247_/A _08018_/B vssd1 vssd1 vccd1 vccd1 _08198_/B sky130_fd_sc_hd__xnor2_2
XFILLER_150_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09969_ _09965_/Y _09968_/X _09894_/X vssd1 vssd1 vccd1 vccd1 _09969_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12980_ _12978_/A _12978_/B _12979_/X vssd1 vssd1 vccd1 vccd1 _16188_/D sky130_fd_sc_hd__a21oi_1
XFILLER_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11931_ _11927_/Y _11928_/X _11930_/Y _11925_/C vssd1 vssd1 vccd1 vccd1 _11933_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_73_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14650_ _14648_/Y _14643_/C _14645_/Y _14646_/X vssd1 vssd1 vccd1 vccd1 _14651_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_45_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11862_ _16032_/Q _11869_/C _11748_/X vssd1 vssd1 vccd1 vccd1 _11865_/B sky130_fd_sc_hd__a21o_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13601_ _13635_/A _13601_/B _13601_/C vssd1 vssd1 vccd1 vccd1 _13602_/A sky130_fd_sc_hd__and3_1
XFILLER_26_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10813_ _10813_/A _10823_/B vssd1 vssd1 vccd1 vccd1 _10816_/A sky130_fd_sc_hd__or2_1
X_14581_ _16420_/Q _14583_/C _14411_/X vssd1 vssd1 vccd1 vccd1 _14581_/Y sky130_fd_sc_hd__a21oi_1
X_11793_ input7/X vssd1 vssd1 vccd1 vccd1 _12924_/A sky130_fd_sc_hd__buf_2
X_16320_ _16346_/CLK _16320_/D vssd1 vssd1 vccd1 vccd1 _16320_/Q sky130_fd_sc_hd__dfxtp_1
X_13532_ _14095_/A vssd1 vssd1 vccd1 vccd1 _13760_/B sky130_fd_sc_hd__clkbuf_2
X_10744_ _10741_/Y _10742_/X _10743_/Y _10738_/C vssd1 vssd1 vccd1 vccd1 _10746_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16251_ _16261_/CLK _16251_/D vssd1 vssd1 vccd1 vccd1 _16251_/Q sky130_fd_sc_hd__dfxtp_1
X_13463_ _13463_/A vssd1 vssd1 vccd1 vccd1 _16257_/D sky130_fd_sc_hd__clkbuf_1
X_10675_ _15861_/Q _10726_/B _10675_/C vssd1 vssd1 vccd1 vccd1 _10681_/A sky130_fd_sc_hd__and3_1
XFILLER_139_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15202_ _16519_/Q _15255_/B _15209_/C vssd1 vssd1 vccd1 vccd1 _15202_/Y sky130_fd_sc_hd__nand3_1
X_12414_ _12412_/A _12412_/B _12413_/X vssd1 vssd1 vccd1 vccd1 _16108_/D sky130_fd_sc_hd__a21oi_1
X_16182_ _16237_/CLK _16182_/D vssd1 vssd1 vccd1 vccd1 _16182_/Q sky130_fd_sc_hd__dfxtp_2
X_13394_ _13391_/Y _13393_/X _13388_/C _13389_/C vssd1 vssd1 vccd1 vccd1 _13396_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_139_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15133_ _15133_/A vssd1 vssd1 vccd1 vccd1 _16507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12345_ _16100_/Q _12352_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12345_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15064_ _15117_/A _15064_/B _15064_/C vssd1 vssd1 vccd1 vccd1 _15065_/C sky130_fd_sc_hd__or3_1
XFILLER_142_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12276_ _16091_/Q _12287_/C _12050_/X vssd1 vssd1 vccd1 vccd1 _12276_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ _14015_/A vssd1 vssd1 vccd1 vccd1 _14015_/X sky130_fd_sc_hd__clkbuf_2
X_11227_ _11264_/A _11227_/B _11227_/C vssd1 vssd1 vccd1 vccd1 _11228_/A sky130_fd_sc_hd__and3_1
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11158_ _12292_/A vssd1 vssd1 vccd1 vccd1 _11158_/X sky130_fd_sc_hd__buf_2
XFILLER_95_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10109_ _10109_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__nor2_1
X_15966_ _16005_/CLK _15966_/D vssd1 vssd1 vccd1 vccd1 _15966_/Q sky130_fd_sc_hd__dfxtp_2
X_11089_ _11089_/A vssd1 vssd1 vccd1 vccd1 _15922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14917_ _16473_/Q _14925_/C _14858_/X vssd1 vssd1 vccd1 vccd1 _14917_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15897_ _16553_/Q _15897_/D vssd1 vssd1 vccd1 vccd1 _15897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16632__37 vssd1 vssd1 vccd1 vccd1 _16632__37/HI _16698_/A sky130_fd_sc_hd__conb_1
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14848_ _14848_/A vssd1 vssd1 vccd1 vccd1 _15074_/B sky130_fd_sc_hd__clkbuf_2
X_14779_ _14780_/B _14780_/C _14669_/X vssd1 vssd1 vccd1 vccd1 _14781_/B sky130_fd_sc_hd__o21ai_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16518_ _16607_/CLK _16518_/D vssd1 vssd1 vccd1 vccd1 _16518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16449_ _16607_/CLK _16449_/D vssd1 vssd1 vccd1 vccd1 _16449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09823_ _13288_/A vssd1 vssd1 vccd1 vccd1 _14979_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09754_ _09617_/X _09706_/X _09747_/B _09707_/X vssd1 vssd1 vccd1 vccd1 _09755_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_86_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08705_ _09038_/A _08705_/B _08705_/C vssd1 vssd1 vccd1 vccd1 _08710_/A sky130_fd_sc_hd__and3_1
XFILLER_104_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09685_ _15255_/B vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ input5/X vssd1 vssd1 vccd1 vccd1 _12849_/A sky130_fd_sc_hd__buf_6
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08567_ _08567_/A _08567_/B vssd1 vssd1 vccd1 vccd1 _08567_/X sky130_fd_sc_hd__or2_1
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08498_ _08459_/A _08459_/B _08461_/B vssd1 vssd1 vccd1 vccd1 _08499_/B sky130_fd_sc_hd__a21oi_1
XFILLER_120_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10460_ _10458_/Y _10451_/C _10455_/Y _10465_/A vssd1 vssd1 vccd1 vccd1 _10465_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_6_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ _09119_/A _09124_/C vssd1 vssd1 vccd1 vccd1 _09119_/Y sky130_fd_sc_hd__nor2_1
X_10391_ _10399_/A _10391_/B _10391_/C vssd1 vssd1 vccd1 vccd1 _10392_/A sky130_fd_sc_hd__and3_1
XFILLER_135_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12130_ _12128_/A _12128_/B _12129_/X vssd1 vssd1 vccd1 vccd1 _16068_/D sky130_fd_sc_hd__a21oi_1
XFILLER_135_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12061_ _12058_/Y _12067_/A _12060_/Y _12056_/C vssd1 vssd1 vccd1 vccd1 _12063_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ _15912_/Q _11183_/B _11018_/C vssd1 vssd1 vccd1 vccd1 _11014_/C sky130_fd_sc_hd__nand3_1
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15820_ _16551_/CLK _15820_/D vssd1 vssd1 vccd1 vccd1 _15820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15751_ _15791_/CLK _15751_/D vssd1 vssd1 vccd1 vccd1 _15751_/Q sky130_fd_sc_hd__dfxtp_2
X_12963_ _12963_/A _12963_/B _12963_/C vssd1 vssd1 vccd1 vccd1 _12964_/A sky130_fd_sc_hd__and3_1
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14702_ _16439_/Q _14710_/C _14588_/X vssd1 vssd1 vccd1 vccd1 _14702_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11914_ _11948_/A _11914_/B _11918_/A vssd1 vssd1 vccd1 vccd1 _16038_/D sky130_fd_sc_hd__nor3_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _15791_/CLK _15682_/D vssd1 vssd1 vccd1 vccd1 _15682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12894_ _16178_/Q _12896_/C _12723_/X vssd1 vssd1 vccd1 vccd1 _12894_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _16428_/Q _14742_/B _14633_/C vssd1 vssd1 vccd1 vccd1 _14633_/X sky130_fd_sc_hd__and3_1
X_11845_ _11845_/A _11845_/B vssd1 vssd1 vccd1 vccd1 _11846_/B sky130_fd_sc_hd__nor2_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14564_ _14848_/A vssd1 vssd1 vccd1 vccd1 _14790_/B sky130_fd_sc_hd__buf_2
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _11776_/A _11776_/B _11776_/C vssd1 vssd1 vccd1 vccd1 _11777_/A sky130_fd_sc_hd__and3_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16533_/Q _16303_/D vssd1 vssd1 vccd1 vccd1 _16303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13515_ _13512_/Y _13513_/X _13514_/Y _13510_/C vssd1 vssd1 vccd1 vccd1 _13517_/B
+ sky130_fd_sc_hd__o211ai_1
X_10727_ _10809_/A _10727_/B _10731_/A vssd1 vssd1 vccd1 vccd1 _15868_/D sky130_fd_sc_hd__nor3_1
X_14495_ _14496_/B _14496_/C _14387_/X vssd1 vssd1 vccd1 vccd1 _14497_/B sky130_fd_sc_hd__o21ai_1
XFILLER_146_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ _16261_/CLK _16234_/D vssd1 vssd1 vccd1 vccd1 _16234_/Q sky130_fd_sc_hd__dfxtp_1
X_13446_ _13447_/B _13447_/C _13447_/A vssd1 vssd1 vccd1 vccd1 _13448_/B sky130_fd_sc_hd__a21o_1
X_10658_ _15857_/Q _10707_/B _10658_/C vssd1 vssd1 vccd1 vccd1 _10659_/B sky130_fd_sc_hd__and3_1
XFILLER_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16165_ _16237_/CLK _16165_/D vssd1 vssd1 vccd1 vccd1 _16165_/Q sky130_fd_sc_hd__dfxtp_1
X_13377_ _13377_/A vssd1 vssd1 vccd1 vccd1 _13498_/A sky130_fd_sc_hd__buf_2
X_10589_ _10589_/A _10589_/B _10589_/C vssd1 vssd1 vccd1 vccd1 _10590_/A sky130_fd_sc_hd__and3_1
X_15116_ _15117_/B _15117_/C _14954_/X vssd1 vssd1 vccd1 vccd1 _15118_/B sky130_fd_sc_hd__o21ai_1
X_12328_ _12343_/A _12328_/B _12328_/C vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__and3_1
XFILLER_127_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16096_ _16118_/CLK _16096_/D vssd1 vssd1 vccd1 vccd1 _16096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15047_ _16494_/Q _15055_/C _14821_/X vssd1 vssd1 vccd1 vccd1 _15047_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12259_ _12259_/A vssd1 vssd1 vccd1 vccd1 _16087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15949_ _15365_/A _15949_/D vssd1 vssd1 vccd1 vccd1 _15949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09470_ _09468_/A _09468_/B _09467_/Y _09469_/Y vssd1 vssd1 vccd1 vccd1 _15628_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08421_ _08109_/C _08309_/Y _08420_/X vssd1 vssd1 vccd1 vccd1 _08421_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08352_ _08169_/A _08169_/B _08350_/X _08351_/Y vssd1 vssd1 vccd1 vccd1 _08353_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08283_ _08283_/A _08283_/B vssd1 vssd1 vccd1 vccd1 _08404_/A sky130_fd_sc_hd__xnor2_4
XFILLER_149_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09806_ _10486_/A vssd1 vssd1 vccd1 vccd1 _10288_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07998_ _11287_/A _07998_/B vssd1 vssd1 vccd1 vccd1 _07999_/B sky130_fd_sc_hd__xnor2_1
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09737_ _09734_/A _09733_/Y _09734_/B vssd1 vssd1 vccd1 vccd1 _09737_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09668_ _15673_/Q _09692_/C _09493_/X vssd1 vssd1 vccd1 vccd1 _09670_/B sky130_fd_sc_hd__a21oi_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _15461_/Q _09271_/A _08619_/C vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__and3_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09599_ _09599_/A _09599_/B vssd1 vssd1 vccd1 vccd1 _09599_/X sky130_fd_sc_hd__or2_1
XFILLER_43_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11666_/A _11630_/B _11634_/A vssd1 vssd1 vccd1 vccd1 _15998_/D sky130_fd_sc_hd__nor3_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ _11561_/A _11569_/B vssd1 vssd1 vccd1 vccd1 _11563_/A sky130_fd_sc_hd__or2_1
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13300_ _13297_/Y _13298_/X _13299_/Y _13295_/C vssd1 vssd1 vccd1 vccd1 _13302_/B
+ sky130_fd_sc_hd__o211ai_1
X_10512_ _10508_/Y _10519_/A _10511_/Y _10506_/C vssd1 vssd1 vccd1 vccd1 _10514_/B
+ sky130_fd_sc_hd__o211a_1
X_14280_ _14296_/C vssd1 vssd1 vccd1 vccd1 _14303_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11492_ _11492_/A vssd1 vssd1 vccd1 vccd1 _15978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13231_ _13246_/A _13231_/B _13231_/C vssd1 vssd1 vccd1 vccd1 _13232_/A sky130_fd_sc_hd__and3_1
XFILLER_10_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10443_ _10497_/A _10443_/B _10443_/C vssd1 vssd1 vccd1 vccd1 _10444_/A sky130_fd_sc_hd__and3_1
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13162_ _13443_/A vssd1 vssd1 vccd1 vccd1 _13162_/X sky130_fd_sc_hd__clkbuf_2
X_10374_ _15794_/Q _15793_/Q _15792_/Q _10227_/X vssd1 vssd1 vccd1 vccd1 _15804_/D
+ sky130_fd_sc_hd__o31a_1
X_12113_ _12113_/A _12113_/B _12113_/C vssd1 vssd1 vccd1 vccd1 _12114_/A sky130_fd_sc_hd__and3_1
XFILLER_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ _13151_/A _13093_/B _13093_/C vssd1 vssd1 vccd1 vccd1 _13094_/C sky130_fd_sc_hd__or3_1
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12044_ _16058_/Q _12210_/B _12045_/C vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__and3_1
XFILLER_78_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15803_ _15812_/CLK _15803_/D vssd1 vssd1 vccd1 vccd1 _15803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13995_ _14160_/A vssd1 vssd1 vccd1 vccd1 _14035_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15734_ _16551_/CLK _15734_/D vssd1 vssd1 vccd1 vccd1 _15734_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12946_ _12944_/Y _12945_/X _12941_/C _12942_/C vssd1 vssd1 vccd1 vccd1 _12948_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15665_ _15791_/CLK _15665_/D vssd1 vssd1 vccd1 vccd1 _15665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12877_ _16175_/Q _13102_/B _12889_/C vssd1 vssd1 vccd1 vccd1 _12883_/A sky130_fd_sc_hd__and3_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _16414_/Q _16413_/Q _16412_/Q _14615_/X vssd1 vssd1 vccd1 vccd1 _16424_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _11828_/A vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__clkbuf_2
X_15596_ _16551_/CLK _15596_/D vssd1 vssd1 vccd1 vccd1 _15596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _16414_/Q _14770_/B _14547_/C vssd1 vssd1 vccd1 vccd1 _14555_/B sky130_fd_sc_hd__and3_1
X_11759_ _11752_/C _11753_/C _11756_/Y _11757_/X vssd1 vssd1 vccd1 vccd1 _11760_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14478_ _16404_/Q _14486_/C _14258_/X vssd1 vssd1 vccd1 vccd1 _14478_/Y sky130_fd_sc_hd__a21oi_1
X_16217_ _16237_/CLK _16217_/D vssd1 vssd1 vccd1 vccd1 _16217_/Q sky130_fd_sc_hd__dfxtp_1
X_13429_ _13427_/A _13427_/B _13428_/X vssd1 vssd1 vccd1 vccd1 _16252_/D sky130_fd_sc_hd__a21oi_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16148_ _16555_/Q _16148_/D vssd1 vssd1 vccd1 vccd1 _16148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08970_ _09400_/A vssd1 vssd1 vccd1 vccd1 _09054_/A sky130_fd_sc_hd__clkbuf_2
X_16079_ _16118_/CLK _16079_/D vssd1 vssd1 vccd1 vccd1 _16079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07921_ _16604_/Q _16602_/Q vssd1 vssd1 vccd1 vccd1 _07922_/B sky130_fd_sc_hd__or2_1
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07852_ _15207_/A vssd1 vssd1 vccd1 vccd1 _15367_/B sky130_fd_sc_hd__buf_4
XFILLER_69_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07783_ _07787_/A vssd1 vssd1 vccd1 vccd1 _07783_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09522_ _09517_/Y _09521_/X _09431_/X vssd1 vssd1 vccd1 vccd1 _09522_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09453_ _09453_/A _09453_/B _09453_/C vssd1 vssd1 vccd1 vccd1 _09454_/C sky130_fd_sc_hd__nand3_1
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08404_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08404_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09384_ _15614_/Q _09382_/C _09383_/X vssd1 vssd1 vccd1 vccd1 _09385_/B sky130_fd_sc_hd__a21o_1
X_08335_ _08336_/A _08336_/B _08336_/C vssd1 vssd1 vccd1 vccd1 _08443_/A sky130_fd_sc_hd__a21o_1
XFILLER_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08266_ _15121_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08266_/X sky130_fd_sc_hd__or2_1
XFILLER_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08197_ _08197_/A vssd1 vssd1 vccd1 vccd1 _08197_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16668__73 vssd1 vssd1 vccd1 vccd1 _16668__73/HI _16744_/A sky130_fd_sc_hd__conb_1
X_10090_ _10090_/A vssd1 vssd1 vccd1 vccd1 _15753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12800_ _12800_/A _12800_/B vssd1 vssd1 vccd1 vccd1 _12802_/B sky130_fd_sc_hd__nor2_1
XFILLER_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13780_ _13815_/C vssd1 vssd1 vccd1 vccd1 _13822_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10992_ _15909_/Q _11099_/B _10992_/C vssd1 vssd1 vccd1 vccd1 _11001_/B sky130_fd_sc_hd__and3_1
XFILLER_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _16155_/Q _12739_/C _12619_/X vssd1 vssd1 vccd1 vccd1 _12731_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _16570_/CLK _15450_/D vssd1 vssd1 vccd1 vccd1 _15450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12662_ _16145_/Q _12670_/C _12605_/X vssd1 vssd1 vccd1 vccd1 _12662_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14402_/B _14402_/C _14402_/A vssd1 vssd1 vccd1 vccd1 _14403_/B sky130_fd_sc_hd__a21o_1
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _15997_/Q _11668_/B _11613_/C vssd1 vssd1 vccd1 vccd1 _11621_/B sky130_fd_sc_hd__and3_1
X_15381_ _15973_/Q _15972_/Q _15971_/Q _15378_/X vssd1 vssd1 vccd1 vccd1 _16567_/D
+ sky130_fd_sc_hd__o31a_1
X_12593_ _16135_/Q _12634_/C _12368_/X vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__a21oi_1
X_14332_ _14555_/A _14332_/B _14332_/C vssd1 vssd1 vccd1 vccd1 _14333_/C sky130_fd_sc_hd__or3_1
X_11544_ _15986_/Q _11773_/B _11551_/C vssd1 vssd1 vccd1 vccd1 _11544_/Y sky130_fd_sc_hd__nand3_1
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14263_ _14261_/Y _14256_/C _14259_/Y _14270_/A vssd1 vssd1 vccd1 vccd1 _14270_/B
+ sky130_fd_sc_hd__a211oi_1
X_11475_ _11467_/C _11468_/C _11472_/Y _11473_/X vssd1 vssd1 vccd1 vccd1 _11476_/C
+ sky130_fd_sc_hd__a211o_1
X_16002_ _16005_/CLK _16002_/D vssd1 vssd1 vccd1 vccd1 _16002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ _13235_/C vssd1 vssd1 vccd1 vccd1 _13250_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10426_ _11233_/A vssd1 vssd1 vccd1 vccd1 _10426_/X sky130_fd_sc_hd__clkbuf_2
X_14194_ _16362_/Q _14311_/B _14201_/C vssd1 vssd1 vccd1 vccd1 _14194_/Y sky130_fd_sc_hd__nand3_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13145_ _13145_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _13146_/B sky130_fd_sc_hd__nor2_1
X_10357_ _10354_/Y _10364_/A _10356_/Y _10352_/C vssd1 vssd1 vccd1 vccd1 _10359_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _16204_/Q _13305_/B _13076_/C vssd1 vssd1 vccd1 vccd1 _13084_/A sky130_fd_sc_hd__and3_1
XFILLER_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10288_ _15790_/Q _10294_/B _10288_/C vssd1 vssd1 vccd1 vccd1 _10290_/C sky130_fd_sc_hd__nand3_1
X_12027_ _16055_/Q _12252_/B _12038_/C vssd1 vssd1 vccd1 vccd1 _12033_/A sky130_fd_sc_hd__and3_1
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13978_ _13978_/A vssd1 vssd1 vccd1 vccd1 _16330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15717_ _15812_/CLK _15717_/D vssd1 vssd1 vccd1 vccd1 _15717_/Q sky130_fd_sc_hd__dfxtp_2
X_12929_ _12945_/C vssd1 vssd1 vccd1 vccd1 _12952_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16697_ _16697_/A _07796_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15648_ _15791_/CLK _15648_/D vssd1 vssd1 vccd1 vccd1 _15648_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15579_ _15812_/CLK _15579_/D vssd1 vssd1 vccd1 vccd1 _15579_/Q sky130_fd_sc_hd__dfxtp_1
X_08120_ _12987_/A _07874_/B _07877_/A vssd1 vssd1 vccd1 vccd1 _08143_/A sky130_fd_sc_hd__o21bai_4
XFILLER_147_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08051_ _08051_/A _08228_/A vssd1 vssd1 vccd1 vccd1 _08200_/B sky130_fd_sc_hd__xor2_4
XFILLER_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08953_ _08951_/A _08951_/B _08952_/X vssd1 vssd1 vccd1 vccd1 _15520_/D sky130_fd_sc_hd__a21oi_1
X_07904_ _16572_/Q vssd1 vssd1 vccd1 vccd1 _11683_/A sky130_fd_sc_hd__inv_2
XFILLER_130_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ _08796_/X _08882_/A _08711_/X vssd1 vssd1 vccd1 vccd1 _08884_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07835_ _07836_/A vssd1 vssd1 vccd1 vccd1 _07835_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07766_ _07768_/A vssd1 vssd1 vccd1 vccd1 _07766_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09505_ _09953_/A vssd1 vssd1 vccd1 vccd1 _09595_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09436_/B vssd1 vssd1 vccd1 vccd1 _09436_/Y sky130_fd_sc_hd__nor2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09367_/A _09367_/B _09367_/C vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__and3_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08318_ _08318_/A _08144_/A vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__or2b_1
XFILLER_138_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09298_ _15358_/B vssd1 vssd1 vccd1 vccd1 _09749_/A sky130_fd_sc_hd__clkbuf_2
X_08249_ _09496_/C _08065_/B _08064_/A vssd1 vssd1 vccd1 vccd1 _08251_/C sky130_fd_sc_hd__o21a_1
X_11260_ _11828_/A vssd1 vssd1 vccd1 vccd1 _11488_/B sky130_fd_sc_hd__buf_2
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10211_ _10311_/A _10211_/B _10216_/B vssd1 vssd1 vccd1 vccd1 _15773_/D sky130_fd_sc_hd__nor3_1
XFILLER_134_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11191_ _11189_/Y _11190_/X _11185_/C _11186_/C vssd1 vssd1 vccd1 vccd1 _11193_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_133_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10142_ _15764_/Q _10396_/B _10152_/C vssd1 vssd1 vccd1 vccd1 _10142_/Y sky130_fd_sc_hd__nand3_1
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ _10086_/C vssd1 vssd1 vccd1 vccd1 _10099_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14950_ _14950_/A _14950_/B vssd1 vssd1 vccd1 vccd1 _14956_/C sky130_fd_sc_hd__nor2_1
XFILLER_121_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13901_ _13899_/Y _13900_/X _13896_/C _13897_/C vssd1 vssd1 vccd1 vccd1 _13903_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14881_ _16467_/Q _14995_/B _14881_/C vssd1 vssd1 vccd1 vccd1 _14889_/A sky130_fd_sc_hd__and3_1
XFILLER_63_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13832_ _13866_/A _13832_/B _13832_/C vssd1 vssd1 vccd1 vccd1 _13833_/A sky130_fd_sc_hd__and3_1
XFILLER_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16551_ _16551_/CLK _16551_/D vssd1 vssd1 vccd1 vccd1 _16551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13763_ _13784_/A _13763_/B _13767_/B vssd1 vssd1 vccd1 vccd1 _16299_/D sky130_fd_sc_hd__nor3_1
X_10975_ _15907_/Q _10985_/C _10919_/X vssd1 vssd1 vccd1 vccd1 _10975_/Y sky130_fd_sc_hd__a21oi_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _12714_/A _12714_/B _12714_/C vssd1 vssd1 vccd1 vccd1 _12715_/C sky130_fd_sc_hd__nand3_1
X_15502_ _16570_/CLK _15502_/D vssd1 vssd1 vccd1 vccd1 _15502_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16482_ _16607_/CLK _16482_/D vssd1 vssd1 vccd1 vccd1 _16482_/Q sky130_fd_sc_hd__dfxtp_1
X_13694_ _13689_/Y _13692_/X _13693_/Y _13687_/C vssd1 vssd1 vccd1 vccd1 _13696_/B
+ sky130_fd_sc_hd__o211ai_1
X_15433_ _16309_/Q _16308_/Q _16307_/Q _15428_/X vssd1 vssd1 vccd1 vccd1 _16609_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12645_ _12645_/A vssd1 vssd1 vccd1 vccd1 _16141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15364_ _16711_/A _16710_/A _16709_/A _15363_/X vssd1 vssd1 vccd1 vccd1 _16552_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12576_ _16133_/Q _12578_/C _12575_/X vssd1 vssd1 vccd1 vccd1 _12579_/A sky130_fd_sc_hd__a21oi_1
X_14315_ _14315_/A vssd1 vssd1 vccd1 vccd1 _16378_/D sky130_fd_sc_hd__clkbuf_1
X_11527_ _11527_/A vssd1 vssd1 vccd1 vccd1 _15983_/D sky130_fd_sc_hd__clkbuf_1
X_15295_ _15292_/X _15294_/X _10716_/X vssd1 vssd1 vccd1 vccd1 _15295_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14246_ _14242_/Y _14244_/X _14245_/Y _14240_/C vssd1 vssd1 vccd1 vccd1 _14248_/B
+ sky130_fd_sc_hd__o211ai_1
X_11458_ _11494_/C vssd1 vssd1 vccd1 vccd1 _11500_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10409_ _10409_/A _10409_/B vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__or2_1
X_14177_ _14177_/A vssd1 vssd1 vccd1 vccd1 _16359_/D sky130_fd_sc_hd__clkbuf_1
X_11389_ _11619_/A vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _16210_/Q _13187_/B _13135_/C vssd1 vssd1 vccd1 vccd1 _13128_/Y sky130_fd_sc_hd__nand3_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _16202_/Q _13059_/B _13062_/C vssd1 vssd1 vccd1 vccd1 _13059_/X sky130_fd_sc_hd__and3_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16749_ _16749_/A _07766_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09221_ _09222_/B _09222_/C _09222_/A vssd1 vssd1 vccd1 vccd1 _09223_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _09152_/A _09152_/B vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__nor2_1
XFILLER_148_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08103_ _08302_/A _08303_/B vssd1 vssd1 vccd1 vccd1 _08104_/B sky130_fd_sc_hd__xnor2_2
X_09083_ _09083_/A _09083_/B vssd1 vssd1 vccd1 vccd1 _15549_/D sky130_fd_sc_hd__nor2_1
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08034_ _08034_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08035_/B sky130_fd_sc_hd__nand2_2
XFILLER_135_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09985_ _09998_/C vssd1 vssd1 vccd1 vccd1 _10009_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16638__43 vssd1 vssd1 vccd1 vccd1 _16638__43/HI _16714_/A sky130_fd_sc_hd__conb_1
XFILLER_103_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08936_ _15522_/Q _08937_/C _08805_/X vssd1 vssd1 vccd1 vccd1 _08939_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08867_ _08867_/A _08867_/B vssd1 vssd1 vccd1 vccd1 _08869_/A sky130_fd_sc_hd__or2_1
XFILLER_123_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07818_ _07818_/A vssd1 vssd1 vccd1 vccd1 _07818_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08798_ _08661_/X _08793_/A _08797_/Y vssd1 vssd1 vccd1 vccd1 _15488_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10760_ _10758_/A _10758_/B _10759_/X vssd1 vssd1 vccd1 vccd1 _15873_/D sky130_fd_sc_hd__a21oi_1
XFILLER_16_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater18 _16533_/Q vssd1 vssd1 vccd1 vccd1 _16346_/CLK sky130_fd_sc_hd__buf_12
X_09419_ _09497_/A _09419_/B _09422_/B vssd1 vssd1 vccd1 vccd1 _15618_/D sky130_fd_sc_hd__nor3_1
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10691_ _15864_/Q _10691_/B _10701_/C vssd1 vssd1 vccd1 vccd1 _10691_/X sky130_fd_sc_hd__and3_1
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12430_ _12431_/B _12431_/C _12431_/A vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12361_ _12586_/A _12361_/B _12361_/C vssd1 vssd1 vccd1 vccd1 _12362_/C sky130_fd_sc_hd__or3_1
X_14100_ _16349_/Q _14101_/C _13986_/X vssd1 vssd1 vccd1 vccd1 _14102_/A sky130_fd_sc_hd__a21oi_1
X_11312_ _11319_/A _11312_/B _11312_/C vssd1 vssd1 vccd1 vccd1 _11313_/A sky130_fd_sc_hd__and3_1
X_15080_ _15100_/A _15080_/B _15080_/C vssd1 vssd1 vccd1 vccd1 _15081_/A sky130_fd_sc_hd__and3_1
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12292_ _12292_/A vssd1 vssd1 vccd1 vccd1 _12292_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14031_ _16339_/Q _14193_/B _14038_/C vssd1 vssd1 vccd1 vccd1 _14031_/X sky130_fd_sc_hd__and3_1
XFILLER_141_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11243_ _11264_/A _11243_/B _11243_/C vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__and3_1
XFILLER_106_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11174_ _11197_/C vssd1 vssd1 vccd1 vccd1 _11211_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10125_ _10179_/A _10125_/B _10129_/A vssd1 vssd1 vccd1 vccd1 _15760_/D sky130_fd_sc_hd__nor3_1
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15982_ _16005_/CLK _15982_/D vssd1 vssd1 vccd1 vccd1 _15982_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10056_ _15749_/Q _10057_/C _09699_/A vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__a21oi_1
X_14933_ _16474_/Q _15149_/B _14940_/C vssd1 vssd1 vccd1 vccd1 _14933_/Y sky130_fd_sc_hd__nand3_1
XFILLER_57_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14864_ _14864_/A vssd1 vssd1 vccd1 vccd1 _16463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _16607_/CLK _16603_/D vssd1 vssd1 vccd1 vccd1 _16603_/Q sky130_fd_sc_hd__dfxtp_1
X_13815_ _16308_/Q _13869_/B _13815_/C vssd1 vssd1 vccd1 vccd1 _13824_/A sky130_fd_sc_hd__and3_1
X_14795_ _14795_/A _14795_/B _14795_/C vssd1 vssd1 vccd1 vccd1 _14796_/C sky130_fd_sc_hd__nand3_1
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16534_ _16607_/CLK _16534_/D vssd1 vssd1 vccd1 vccd1 _16534_/Q sky130_fd_sc_hd__dfxtp_2
X_13746_ _13743_/Y _13744_/X _13745_/Y _13741_/C vssd1 vssd1 vccd1 vccd1 _13748_/B
+ sky130_fd_sc_hd__o211ai_1
X_10958_ _10959_/B _10959_/C _10959_/A vssd1 vssd1 vccd1 vccd1 _10960_/B sky130_fd_sc_hd__a21o_1
X_13677_ _13673_/Y _13676_/X _13670_/C _13671_/C vssd1 vssd1 vccd1 vccd1 _13679_/B
+ sky130_fd_sc_hd__o211ai_1
X_16465_ _16607_/CLK _16465_/D vssd1 vssd1 vccd1 vccd1 _16465_/Q sky130_fd_sc_hd__dfxtp_1
X_10889_ _10889_/A vssd1 vssd1 vccd1 vccd1 _10907_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15416_ _15440_/A vssd1 vssd1 vccd1 vccd1 _15416_/X sky130_fd_sc_hd__clkbuf_4
X_12628_ _16140_/Q _12739_/B _12628_/C vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__and3_1
X_16396_ input11/X _16396_/D vssd1 vssd1 vccd1 vccd1 _16396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15347_ _15347_/A _15347_/B vssd1 vssd1 vccd1 vccd1 _15349_/A sky130_fd_sc_hd__or2_1
XFILLER_129_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12559_ _16131_/Q _12569_/C _12337_/X vssd1 vssd1 vccd1 vccd1 _12559_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15278_ _16533_/Q _15366_/B vssd1 vssd1 vccd1 vccd1 _16533_/D sky130_fd_sc_hd__nor2_1
X_14229_ _16368_/Q _14237_/C _14008_/X vssd1 vssd1 vccd1 vccd1 _14232_/B sky130_fd_sc_hd__a21o_1
XFILLER_132_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ _15693_/Q _09914_/B _09770_/C vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__and3_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _15477_/Q _08807_/B _08721_/C vssd1 vssd1 vccd1 vccd1 _08723_/C sky130_fd_sc_hd__nand3_1
XFILLER_79_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08652_ _09164_/A vssd1 vssd1 vccd1 vccd1 _09898_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_39_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08583_ _10486_/A vssd1 vssd1 vccd1 vccd1 _09056_/A sky130_fd_sc_hd__buf_2
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09204_ _15358_/A _15358_/B _09204_/C vssd1 vssd1 vccd1 vccd1 _09206_/A sky130_fd_sc_hd__and3_1
XFILLER_10_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09135_ _15566_/Q _09150_/C _09051_/X vssd1 vssd1 vccd1 vccd1 _09137_/B sky130_fd_sc_hd__a21oi_1
XFILLER_148_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09066_ _09064_/Y _09072_/A _09059_/C _09060_/C vssd1 vssd1 vccd1 vccd1 _09068_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08017_ _12364_/A _08222_/B vssd1 vssd1 vccd1 vccd1 _08018_/B sky130_fd_sc_hd__xnor2_1
XFILLER_118_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09968_ _09966_/X _09968_/B vssd1 vssd1 vccd1 vccd1 _09968_/X sky130_fd_sc_hd__and2b_1
XFILLER_58_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08919_ _08832_/X _08921_/C _08833_/X vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__o21ai_1
X_09899_ _10220_/A _09706_/X _09891_/B _09707_/X vssd1 vssd1 vccd1 vccd1 _09900_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11930_ _16041_/Q _12160_/B _11930_/C vssd1 vssd1 vccd1 vccd1 _11930_/Y sky130_fd_sc_hd__nand3_1
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ _11948_/A _11861_/B _11865_/A vssd1 vssd1 vccd1 vccd1 _16030_/D sky130_fd_sc_hd__nor3_1
XFILLER_73_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13600_ _13717_/A _13600_/B _13600_/C vssd1 vssd1 vccd1 vccd1 _13601_/C sky130_fd_sc_hd__or3_1
X_10812_ _15884_/Q _10812_/B _10812_/C vssd1 vssd1 vccd1 vccd1 _10823_/B sky130_fd_sc_hd__and3_1
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14580_ _14580_/A vssd1 vssd1 vccd1 vccd1 _16418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11792_ _11795_/B _11795_/C _11567_/X vssd1 vssd1 vccd1 vccd1 _11796_/B sky130_fd_sc_hd__o21ai_1
X_13531_ _16268_/Q _13586_/B _13531_/C vssd1 vssd1 vccd1 vccd1 _13540_/A sky130_fd_sc_hd__and3_1
X_10743_ _15872_/Q _10743_/B _10749_/C vssd1 vssd1 vccd1 vccd1 _10743_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ _16261_/CLK _16250_/D vssd1 vssd1 vccd1 vccd1 _16250_/Q sky130_fd_sc_hd__dfxtp_1
X_13462_ _13470_/A _13462_/B _13462_/C vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__and3_1
X_10674_ _15861_/Q _10707_/C _10673_/X vssd1 vssd1 vccd1 vccd1 _10676_/B sky130_fd_sc_hd__a21oi_1
X_15201_ _16520_/Q _15254_/B _15209_/C vssd1 vssd1 vccd1 vccd1 _15201_/X sky130_fd_sc_hd__and3_1
X_12413_ _12466_/A _12418_/C vssd1 vssd1 vccd1 vccd1 _12413_/X sky130_fd_sc_hd__or2_1
X_16181_ _16555_/Q _16181_/D vssd1 vssd1 vccd1 vccd1 _16181_/Q sky130_fd_sc_hd__dfxtp_1
X_13393_ _16249_/Q _13617_/B _13393_/C vssd1 vssd1 vccd1 vccd1 _13393_/X sky130_fd_sc_hd__and3_1
X_15132_ _15152_/A _15132_/B _15132_/C vssd1 vssd1 vccd1 vccd1 _15133_/A sky130_fd_sc_hd__and3_1
XFILLER_127_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12344_ _12344_/A vssd1 vssd1 vccd1 vccd1 _16098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ _15064_/B _15064_/C _14954_/X vssd1 vssd1 vccd1 vccd1 _15065_/B sky130_fd_sc_hd__o21ai_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12275_ _12275_/A vssd1 vssd1 vccd1 vccd1 _16089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14014_ _14014_/A vssd1 vssd1 vccd1 vccd1 _16335_/D sky130_fd_sc_hd__clkbuf_1
X_11226_ _11452_/A _11226_/B _11226_/C vssd1 vssd1 vccd1 vccd1 _11227_/C sky130_fd_sc_hd__or3_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11157_ _12574_/A vssd1 vssd1 vccd1 vccd1 _12292_/A sky130_fd_sc_hd__clkbuf_4
X_10108_ _10108_/A _10108_/B vssd1 vssd1 vccd1 vccd1 _10109_/B sky130_fd_sc_hd__nor2_1
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15965_ _16005_/CLK _15965_/D vssd1 vssd1 vccd1 vccd1 _15965_/Q sky130_fd_sc_hd__dfxtp_1
X_11088_ _11088_/A _11088_/B _11088_/C vssd1 vssd1 vccd1 vccd1 _11089_/A sky130_fd_sc_hd__and3_1
XFILLER_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10039_ _10037_/Y _10038_/X _10034_/C _10035_/C vssd1 vssd1 vccd1 vccd1 _10041_/B
+ sky130_fd_sc_hd__o211ai_1
X_14916_ _14916_/A vssd1 vssd1 vccd1 vccd1 _16471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15896_ _16553_/Q _15896_/D vssd1 vssd1 vccd1 vccd1 _15896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14847_ _16462_/Q _14887_/C _14621_/X vssd1 vssd1 vccd1 vccd1 _14850_/B sky130_fd_sc_hd__a21oi_1
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14778_ _15007_/A vssd1 vssd1 vccd1 vccd1 _14819_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16517_ _16595_/CLK _16517_/D vssd1 vssd1 vccd1 vccd1 _16517_/Q sky130_fd_sc_hd__dfxtp_1
X_13729_ _14851_/A vssd1 vssd1 vccd1 vccd1 _13729_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16448_ _16607_/CLK _16448_/D vssd1 vssd1 vccd1 vccd1 _16448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16379_ _16389_/CLK _16379_/D vssd1 vssd1 vccd1 vccd1 _16379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09822_ _15702_/Q _09836_/C _10003_/B vssd1 vssd1 vccd1 vccd1 _09822_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09753_ _09615_/X _09747_/B _09572_/X vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__a21oi_1
XFILLER_101_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08704_ _08704_/A _08704_/B vssd1 vssd1 vccd1 vccd1 _15468_/D sky130_fd_sc_hd__nor2_1
XFILLER_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09684_ _15676_/Q _09692_/C _09683_/X vssd1 vssd1 vccd1 vccd1 _09688_/A sky130_fd_sc_hd__a21oi_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08635_ _08630_/X _08620_/B _08623_/B _08634_/Y vssd1 vssd1 vccd1 vccd1 _15458_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08566_ _15366_/B _08566_/B _08565_/X vssd1 vssd1 vccd1 vccd1 _15452_/D sky130_fd_sc_hd__nor3b_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08497_ _08497_/A _08497_/B vssd1 vssd1 vccd1 vccd1 _08538_/A sky130_fd_sc_hd__or2_1
XFILLER_120_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09118_ _09111_/B _09115_/B _09117_/X vssd1 vssd1 vccd1 vccd1 _09124_/C sky130_fd_sc_hd__o21a_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10390_ _10384_/C _10385_/C _10387_/Y _10388_/X vssd1 vssd1 vccd1 vccd1 _10391_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ _09057_/C vssd1 vssd1 vccd1 vccd1 _09070_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12060_ _16059_/Q _12060_/B _12065_/C vssd1 vssd1 vccd1 vccd1 _12060_/Y sky130_fd_sc_hd__nand3_1
XFILLER_150_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11011_ _15912_/Q _11018_/C _10898_/X vssd1 vssd1 vccd1 vccd1 _11014_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15750_ _15812_/CLK _15750_/D vssd1 vssd1 vccd1 vccd1 _15750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12962_ _12960_/Y _12955_/C _12957_/Y _12958_/X vssd1 vssd1 vccd1 vccd1 _12963_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14701_ _14701_/A vssd1 vssd1 vccd1 vccd1 _16437_/D sky130_fd_sc_hd__clkbuf_1
X_11913_ _16039_/Q _11969_/B _11922_/C vssd1 vssd1 vccd1 vccd1 _11918_/A sky130_fd_sc_hd__and3_1
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _15791_/CLK _15681_/D vssd1 vssd1 vccd1 vccd1 _15681_/Q sky130_fd_sc_hd__dfxtp_2
X_12893_ _12893_/A vssd1 vssd1 vccd1 vccd1 _16176_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11844_ _11844_/A _11852_/B vssd1 vssd1 vccd1 vccd1 _11846_/A sky130_fd_sc_hd__or2_1
X_14632_ _16428_/Q _14640_/C _14574_/X vssd1 vssd1 vccd1 vccd1 _14632_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14563_ _16417_/Q _14603_/C _14339_/X vssd1 vssd1 vccd1 vccd1 _14566_/B sky130_fd_sc_hd__a21oi_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11773_/Y _11767_/C _11771_/Y _11772_/X vssd1 vssd1 vccd1 vccd1 _11776_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16533_/Q _16302_/D vssd1 vssd1 vccd1 vccd1 _16302_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _15870_/Q _10726_/B _10726_/C vssd1 vssd1 vccd1 vccd1 _10731_/A sky130_fd_sc_hd__and3_1
X_13514_ _16265_/Q _13573_/B _13514_/C vssd1 vssd1 vccd1 vccd1 _13514_/Y sky130_fd_sc_hd__nand3_1
X_14494_ _14722_/A vssd1 vssd1 vccd1 vccd1 _14535_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ _16256_/Q _13445_/B _13452_/C vssd1 vssd1 vccd1 vccd1 _13447_/C sky130_fd_sc_hd__nand3_1
X_16233_ _16261_/CLK _16233_/D vssd1 vssd1 vccd1 vccd1 _16233_/Q sky130_fd_sc_hd__dfxtp_1
X_10657_ _15857_/Q _10658_/C _08748_/A vssd1 vssd1 vccd1 vccd1 _10659_/A sky130_fd_sc_hd__a21oi_1
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ _13376_/A vssd1 vssd1 vccd1 vccd1 _16245_/D sky130_fd_sc_hd__clkbuf_1
X_16164_ _16237_/CLK _16164_/D vssd1 vssd1 vccd1 vccd1 _16164_/Q sky130_fd_sc_hd__dfxtp_1
X_10588_ _10588_/A _10588_/B _10588_/C vssd1 vssd1 vccd1 vccd1 _10589_/C sky130_fd_sc_hd__nand3_1
XFILLER_126_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15115_ _15221_/A vssd1 vssd1 vccd1 vccd1 _15152_/A sky130_fd_sc_hd__clkbuf_2
X_12327_ _12320_/C _12321_/C _12324_/Y _12325_/X vssd1 vssd1 vccd1 vccd1 _12328_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16095_ _16118_/CLK _16095_/D vssd1 vssd1 vccd1 vccd1 _16095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15046_ _15046_/A vssd1 vssd1 vccd1 vccd1 _16492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12258_ _12283_/A _12258_/B _12258_/C vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__and3_1
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11209_ _11209_/A vssd1 vssd1 vccd1 vccd1 _15938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ _12189_/A vssd1 vssd1 vccd1 vccd1 _16077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15948_ _15365_/A _15948_/D vssd1 vssd1 vccd1 vccd1 _15948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15879_ _16553_/Q _15879_/D vssd1 vssd1 vccd1 vccd1 _15879_/Q sky130_fd_sc_hd__dfxtp_1
X_08420_ _15448_/Q _08490_/A _15293_/C vssd1 vssd1 vccd1 vccd1 _08420_/X sky130_fd_sc_hd__and3_1
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08351_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08282_ _08400_/A _08400_/B vssd1 vssd1 vccd1 vccd1 _08283_/B sky130_fd_sc_hd__xor2_4
XFILLER_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09805_ _15700_/Q _09816_/C _10729_/B vssd1 vssd1 vccd1 vccd1 _09809_/B sky130_fd_sc_hd__a21o_1
XFILLER_101_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07997_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _07998_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09736_ _09734_/A _09734_/B _09733_/Y _09735_/Y vssd1 vssd1 vccd1 vccd1 _15682_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_28_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09667_ _09679_/C vssd1 vssd1 vccd1 vccd1 _09692_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08618_ _10501_/A vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09598_ _09598_/A _09598_/B vssd1 vssd1 vccd1 vccd1 _09598_/Y sky130_fd_sc_hd__nor2_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08529_/A _08529_/B _08564_/A vssd1 vssd1 vccd1 vccd1 _08549_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11560_ _15989_/Q _11668_/B _11560_/C vssd1 vssd1 vccd1 vccd1 _11569_/B sky130_fd_sc_hd__and3_1
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10511_ _15828_/Q _10702_/B _10517_/C vssd1 vssd1 vccd1 vccd1 _10511_/Y sky130_fd_sc_hd__nand3_1
XFILLER_128_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11491_ _11491_/A _11491_/B _11491_/C vssd1 vssd1 vccd1 vccd1 _11492_/A sky130_fd_sc_hd__and3_1
X_13230_ _13224_/C _13225_/C _13227_/Y _13228_/X vssd1 vssd1 vccd1 vccd1 _13231_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ _10436_/C _10437_/C _10439_/Y _10440_/X vssd1 vssd1 vccd1 vccd1 _10443_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_109_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13161_ _13219_/A _13161_/B _13166_/A vssd1 vssd1 vccd1 vccd1 _16214_/D sky130_fd_sc_hd__nor3_1
X_10373_ _10276_/X _10370_/B _10372_/Y vssd1 vssd1 vccd1 vccd1 _15803_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12112_ _12110_/Y _12103_/C _12105_/Y _12106_/X vssd1 vssd1 vccd1 vccd1 _12113_/C
+ sky130_fd_sc_hd__a211o_1
X_13092_ _13093_/B _13093_/C _12982_/X vssd1 vssd1 vccd1 vccd1 _13094_/B sky130_fd_sc_hd__o21ai_1
XFILLER_123_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12043_ _16058_/Q _12045_/C _11875_/X vssd1 vssd1 vccd1 vccd1 _12043_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_120_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15802_ _15812_/CLK _15802_/D vssd1 vssd1 vccd1 vccd1 _15802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13994_ _13992_/A _13992_/B _13993_/X vssd1 vssd1 vccd1 vccd1 _16332_/D sky130_fd_sc_hd__a21oi_1
XFILLER_105_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15733_ _16551_/CLK _15733_/D vssd1 vssd1 vccd1 vccd1 _15733_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12945_ _16185_/Q _13053_/B _12945_/C vssd1 vssd1 vccd1 vccd1 _12945_/X sky130_fd_sc_hd__and3_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15664_ _15791_/CLK _15664_/D vssd1 vssd1 vccd1 vccd1 _15664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _13725_/A vssd1 vssd1 vccd1 vccd1 _13102_/B sky130_fd_sc_hd__clkbuf_4
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14615_ _14615_/A vssd1 vssd1 vccd1 vccd1 _14615_/X sky130_fd_sc_hd__buf_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _16027_/Q _11936_/B _11836_/C vssd1 vssd1 vccd1 vccd1 _11827_/X sky130_fd_sc_hd__and3_1
X_15595_ _16551_/CLK _15595_/D vssd1 vssd1 vccd1 vccd1 _15595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11756_/Y _11757_/X _11752_/C _11753_/C vssd1 vssd1 vccd1 vccd1 _11760_/B
+ sky130_fd_sc_hd__o211ai_1
X_14546_ _14830_/A vssd1 vssd1 vccd1 vccd1 _14770_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10709_ _10709_/A _10709_/B vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__nor2_1
X_11689_ _11805_/A _11689_/B _11693_/A vssd1 vssd1 vccd1 vccd1 _16006_/D sky130_fd_sc_hd__nor3_1
X_14477_ _14477_/A vssd1 vssd1 vccd1 vccd1 _16402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16216_ _16237_/CLK _16216_/D vssd1 vssd1 vccd1 vccd1 _16216_/Q sky130_fd_sc_hd__dfxtp_1
X_13428_ _13596_/A _13432_/C vssd1 vssd1 vccd1 vccd1 _13428_/X sky130_fd_sc_hd__or2_1
XFILLER_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13359_ _16243_/Q _13474_/B _13364_/C vssd1 vssd1 vccd1 vccd1 _13359_/Y sky130_fd_sc_hd__nand3_1
X_16147_ _16555_/Q _16147_/D vssd1 vssd1 vccd1 vccd1 _16147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16078_ _16118_/CLK _16078_/D vssd1 vssd1 vccd1 vccd1 _16078_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_130_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07920_ _16604_/Q _16602_/Q vssd1 vssd1 vccd1 vccd1 _07922_/A sky130_fd_sc_hd__nand2_1
X_15029_ _15023_/C _15024_/C _15026_/Y _15027_/X vssd1 vssd1 vccd1 vccd1 _15030_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07851_ _09278_/A vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__buf_4
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_6
X_07782_ _07806_/A vssd1 vssd1 vccd1 vccd1 _07787_/A sky130_fd_sc_hd__buf_12
XFILLER_84_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ _09519_/X _09521_/B vssd1 vssd1 vccd1 vccd1 _09521_/X sky130_fd_sc_hd__and2b_1
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09452_ _09453_/B _09453_/C _09453_/A vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__a21o_1
XFILLER_92_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08403_ _08403_/A _08403_/B vssd1 vssd1 vccd1 vccd1 _08473_/A sky130_fd_sc_hd__xnor2_4
XFILLER_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09383_ _09604_/A vssd1 vssd1 vccd1 vccd1 _09383_/X sky130_fd_sc_hd__buf_2
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08334_ _08135_/A _08135_/B _08333_/Y vssd1 vssd1 vccd1 vccd1 _08336_/C sky130_fd_sc_hd__a21oi_1
X_08265_ _08265_/A _08385_/C vssd1 vssd1 vccd1 vccd1 _08268_/A sky130_fd_sc_hd__xnor2_1
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08196_ _08196_/A _08323_/A vssd1 vssd1 vccd1 vccd1 _08287_/A sky130_fd_sc_hd__xnor2_1
XFILLER_118_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16683__88 vssd1 vssd1 vccd1 vccd1 _16683__88/HI _16759_/A sky130_fd_sc_hd__conb_1
XFILLER_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09719_ _15683_/Q _09727_/C _09583_/X vssd1 vssd1 vccd1 vccd1 _09722_/B sky130_fd_sc_hd__a21o_1
X_10991_ _15909_/Q _10992_/C _10874_/X vssd1 vssd1 vccd1 vccd1 _10993_/A sky130_fd_sc_hd__a21oi_1
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12730_ _12730_/A vssd1 vssd1 vccd1 vccd1 _16153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12661_/A vssd1 vssd1 vccd1 vccd1 _16143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _15997_/Q _11613_/C _11441_/X vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__a21oi_1
X_14400_ _16392_/Q _14569_/B _14406_/C vssd1 vssd1 vccd1 vccd1 _14402_/C sky130_fd_sc_hd__nand3_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12628_/C vssd1 vssd1 vccd1 vccd1 _12634_/C sky130_fd_sc_hd__clkbuf_2
X_15380_ _15965_/Q _15964_/Q _15963_/Q _15378_/X vssd1 vssd1 vccd1 vccd1 _16566_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11543_ _11828_/A vssd1 vssd1 vccd1 vccd1 _11773_/B sky130_fd_sc_hd__clkbuf_2
X_14331_ _14331_/A vssd1 vssd1 vccd1 vccd1 _14555_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14262_ _14259_/Y _14270_/A _14261_/Y _14256_/C vssd1 vssd1 vccd1 vccd1 _14264_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11474_ _11472_/Y _11473_/X _11467_/C _11468_/C vssd1 vssd1 vccd1 vccd1 _11476_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_137_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16001_ _16005_/CLK _16001_/D vssd1 vssd1 vccd1 vccd1 _16001_/Q sky130_fd_sc_hd__dfxtp_1
X_13213_ _13228_/C vssd1 vssd1 vccd1 vccd1 _13235_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10425_ _10457_/C vssd1 vssd1 vccd1 vccd1 _10463_/C sky130_fd_sc_hd__clkbuf_2
X_14193_ _16363_/Q _14193_/B _14201_/C vssd1 vssd1 vccd1 vccd1 _14193_/X sky130_fd_sc_hd__and3_1
X_13144_ _13144_/A _13151_/B vssd1 vssd1 vccd1 vccd1 _13146_/A sky130_fd_sc_hd__or2_1
X_10356_ _15801_/Q _10458_/B _10362_/C vssd1 vssd1 vccd1 vccd1 _10356_/Y sky130_fd_sc_hd__nand3_1
XFILLER_124_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13075_ _13638_/A vssd1 vssd1 vccd1 vccd1 _13305_/B sky130_fd_sc_hd__clkbuf_2
X_10287_ _15790_/Q _10294_/B _10181_/X vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__a21o_1
XFILLER_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12026_ _12312_/A vssd1 vssd1 vccd1 vccd1 _12252_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13977_ _13977_/A _13977_/B _13977_/C vssd1 vssd1 vccd1 vccd1 _13978_/A sky130_fd_sc_hd__and3_1
XFILLER_74_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15716_ _15812_/CLK _15716_/D vssd1 vssd1 vccd1 vccd1 _15716_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _12928_/A vssd1 vssd1 vccd1 vccd1 _12945_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16696_ _16696_/A _07795_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15647_ _15791_/CLK _15647_/D vssd1 vssd1 vccd1 vccd1 _15647_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12859_ _13423_/A vssd1 vssd1 vccd1 vccd1 _13082_/B sky130_fd_sc_hd__buf_2
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15578_ _16551_/CLK _15578_/D vssd1 vssd1 vccd1 vccd1 _15578_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14529_ _16412_/Q _14539_/C _14308_/X vssd1 vssd1 vccd1 vccd1 _14529_/Y sky130_fd_sc_hd__a21oi_1
X_08050_ _12473_/A _08229_/B vssd1 vssd1 vccd1 vccd1 _08228_/A sky130_fd_sc_hd__xnor2_4
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08952_ _09074_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _08952_/X sky130_fd_sc_hd__or2_1
XFILLER_103_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07903_ _16570_/Q vssd1 vssd1 vccd1 vccd1 _11572_/A sky130_fd_sc_hd__inv_2
X_08883_ _10276_/A vssd1 vssd1 vccd1 vccd1 _08883_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07834_ _07836_/A vssd1 vssd1 vccd1 vccd1 _07834_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07765_ _07768_/A vssd1 vssd1 vccd1 vccd1 _07765_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _10697_/A vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__clkbuf_4
X_09435_ _15355_/A _09435_/B vssd1 vssd1 vccd1 vccd1 _09436_/B sky130_fd_sc_hd__and2_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ _09366_/A _09366_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09367_/C sky130_fd_sc_hd__nand3_1
X_08317_ _08294_/A _08294_/B _08300_/A vssd1 vssd1 vccd1 vccd1 _08430_/A sky130_fd_sc_hd__o21ai_2
X_09297_ _09291_/X _09295_/B _09296_/Y vssd1 vssd1 vccd1 vccd1 _15594_/D sky130_fd_sc_hd__o21a_1
XANTENNA_40 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08248_ _14902_/A _08248_/B vssd1 vssd1 vccd1 vccd1 _08251_/B sky130_fd_sc_hd__or2_1
XFILLER_119_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08179_ _11908_/A _07968_/B _08178_/Y vssd1 vssd1 vccd1 vccd1 _08190_/A sky130_fd_sc_hd__o21ai_4
XFILLER_119_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10210_ _10208_/Y _10201_/C _10205_/Y _10216_/A vssd1 vssd1 vccd1 vccd1 _10216_/B
+ sky130_fd_sc_hd__a211oi_1
X_11190_ _15937_/Q _11353_/B _11190_/C vssd1 vssd1 vccd1 vccd1 _11190_/X sky130_fd_sc_hd__and3_1
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10141_ _10447_/A vssd1 vssd1 vccd1 vccd1 _10396_/B sky130_fd_sc_hd__buf_2
XFILLER_0_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10072_ _10076_/C vssd1 vssd1 vccd1 vccd1 _10086_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13900_ _16321_/Q _13900_/B _13900_/C vssd1 vssd1 vccd1 vccd1 _13900_/X sky130_fd_sc_hd__and3_1
XFILLER_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14880_ _16467_/Q _14887_/C _14821_/X vssd1 vssd1 vccd1 vccd1 _14880_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13831_ _13997_/A _13831_/B _13831_/C vssd1 vssd1 vccd1 vccd1 _13832_/C sky130_fd_sc_hd__or3_1
XFILLER_90_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16550_ _16551_/CLK _16550_/D vssd1 vssd1 vccd1 vccd1 _16550_/Q sky130_fd_sc_hd__dfxtp_1
X_10974_ _10974_/A vssd1 vssd1 vccd1 vccd1 _15905_/D sky130_fd_sc_hd__clkbuf_1
X_13762_ _13760_/Y _13756_/C _13758_/Y _13767_/A vssd1 vssd1 vccd1 vccd1 _13767_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15501_ _16551_/CLK _15501_/D vssd1 vssd1 vccd1 vccd1 _15501_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ _12714_/B _12714_/C _12714_/A vssd1 vssd1 vccd1 vccd1 _12715_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16481_ _16607_/CLK _16481_/D vssd1 vssd1 vccd1 vccd1 _16481_/Q sky130_fd_sc_hd__dfxtp_1
X_13693_ _16290_/Q _13753_/B _13700_/C vssd1 vssd1 vccd1 vccd1 _13693_/Y sky130_fd_sc_hd__nand3_1
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15432_ _16301_/Q _16300_/Q _16299_/Q _15428_/X vssd1 vssd1 vccd1 vccd1 _16608_/D
+ sky130_fd_sc_hd__o31a_1
X_12644_ _12681_/A _12644_/B _12644_/C vssd1 vssd1 vccd1 vccd1 _12645_/A sky130_fd_sc_hd__and3_1
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15363_ _15378_/A vssd1 vssd1 vccd1 vccd1 _15363_/X sky130_fd_sc_hd__buf_2
XFILLER_62_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12575_ _13705_/A vssd1 vssd1 vccd1 vccd1 _12575_/X sky130_fd_sc_hd__buf_2
X_14314_ _14314_/A _14314_/B _14314_/C vssd1 vssd1 vccd1 vccd1 _14315_/A sky130_fd_sc_hd__and3_1
X_11526_ _11547_/A _11526_/B _11526_/C vssd1 vssd1 vccd1 vccd1 _11527_/A sky130_fd_sc_hd__and3_1
X_15294_ _15283_/C _15286_/Y _15293_/X vssd1 vssd1 vccd1 vccd1 _15294_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11457_ _11480_/C vssd1 vssd1 vccd1 vccd1 _11494_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14245_ _16369_/Q _14414_/B _14245_/C vssd1 vssd1 vccd1 vccd1 _14245_/Y sky130_fd_sc_hd__nand3_1
XFILLER_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10408_ _15812_/Q _10463_/B _10408_/C vssd1 vssd1 vccd1 vccd1 _10409_/B sky130_fd_sc_hd__and3_1
X_14176_ _14197_/A _14176_/B _14176_/C vssd1 vssd1 vccd1 vccd1 _14177_/A sky130_fd_sc_hd__and3_1
X_11388_ _11957_/A vssd1 vssd1 vccd1 vccd1 _11619_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _10339_/A vssd1 vssd1 vccd1 vccd1 _15797_/D sky130_fd_sc_hd__clkbuf_1
X_13127_ _16211_/Q _13350_/B _13135_/C vssd1 vssd1 vccd1 vccd1 _13127_/X sky130_fd_sc_hd__and3_1
XFILLER_140_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _16202_/Q _13062_/C _13006_/X vssd1 vssd1 vccd1 vccd1 _13058_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12009_ _12009_/A vssd1 vssd1 vccd1 vccd1 _12232_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16748_ _16748_/A _07765_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _15585_/Q _09220_/B _09220_/C vssd1 vssd1 vccd1 vccd1 _09222_/C sky130_fd_sc_hd__nand3_1
X_09151_ _09151_/A _09151_/B vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__or2_1
XFILLER_147_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08102_ _08113_/A _08102_/B vssd1 vssd1 vccd1 vccd1 _08303_/B sky130_fd_sc_hd__xnor2_1
X_09082_ _09038_/X _09084_/C _09039_/X vssd1 vssd1 vccd1 vccd1 _09083_/B sky130_fd_sc_hd__o21ai_1
XFILLER_147_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08033_ _15795_/Q _15777_/Q vssd1 vssd1 vccd1 vccd1 _08034_/B sky130_fd_sc_hd__or2_1
XFILLER_143_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09984_ _09987_/C vssd1 vssd1 vccd1 vccd1 _09998_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_115_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08935_ _08946_/A _08935_/B _08939_/A vssd1 vssd1 vccd1 vccd1 _15517_/D sky130_fd_sc_hd__nor3_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08866_ _15506_/Q _08991_/B _08866_/C vssd1 vssd1 vccd1 vccd1 _08867_/B sky130_fd_sc_hd__and3_1
XFILLER_84_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07817_ _07818_/A vssd1 vssd1 vccd1 vccd1 _07817_/Y sky130_fd_sc_hd__inv_2
X_16653__58 vssd1 vssd1 vccd1 vccd1 _16653__58/HI _16729_/A sky130_fd_sc_hd__conb_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08797_ _08796_/X _08793_/A _08711_/X vssd1 vssd1 vccd1 vccd1 _08797_/Y sky130_fd_sc_hd__a21oi_1
Xrepeater19 _16570_/CLK vssd1 vssd1 vccd1 vccd1 _16551_/CLK sky130_fd_sc_hd__buf_12
X_09418_ _09412_/C _09413_/C _09415_/Y _09422_/A vssd1 vssd1 vccd1 vccd1 _09422_/B
+ sky130_fd_sc_hd__a211oi_1
X_10690_ _15864_/Q _10701_/C _09683_/A vssd1 vssd1 vccd1 vccd1 _10690_/Y sky130_fd_sc_hd__a21oi_1
X_09349_ _09301_/X _09347_/B _09304_/X vssd1 vssd1 vccd1 vccd1 _09349_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12360_ _12924_/A vssd1 vssd1 vccd1 vccd1 _12586_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ _11309_/Y _11304_/C _11307_/Y _11308_/X vssd1 vssd1 vccd1 vccd1 _11312_/C
+ sky130_fd_sc_hd__a211o_1
X_12291_ _12371_/A _12291_/B _12298_/B vssd1 vssd1 vccd1 vccd1 _16091_/D sky130_fd_sc_hd__nor3_1
XFILLER_126_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14030_ _16339_/Q _14038_/C _14029_/X vssd1 vssd1 vccd1 vccd1 _14030_/Y sky130_fd_sc_hd__a21oi_1
X_11242_ _11242_/A _11242_/B _11242_/C vssd1 vssd1 vccd1 vccd1 _11243_/C sky130_fd_sc_hd__nand3_1
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11173_ _11190_/C vssd1 vssd1 vccd1 vccd1 _11197_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10124_ _15762_/Q _10178_/B _10124_/C vssd1 vssd1 vccd1 vccd1 _10129_/A sky130_fd_sc_hd__and3_1
XFILLER_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15981_ _16005_/CLK _15981_/D vssd1 vssd1 vccd1 vccd1 _15981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10055_ _10055_/A _10055_/B _10059_/B vssd1 vssd1 vccd1 vccd1 _15746_/D sky130_fd_sc_hd__nor3_1
XFILLER_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14932_ _14932_/A vssd1 vssd1 vccd1 vccd1 _15149_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14863_ _14878_/A _14863_/B _14863_/C vssd1 vssd1 vccd1 vccd1 _14864_/A sky130_fd_sc_hd__and3_1
XFILLER_63_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16602_ _16607_/CLK _16602_/D vssd1 vssd1 vccd1 vccd1 _16602_/Q sky130_fd_sc_hd__dfxtp_1
X_13814_ _16308_/Q _13822_/C _13698_/X vssd1 vssd1 vccd1 vccd1 _13814_/Y sky130_fd_sc_hd__a21oi_1
X_14794_ _14795_/B _14795_/C _14795_/A vssd1 vssd1 vccd1 vccd1 _14796_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16533_ _16607_/CLK _16533_/D vssd1 vssd1 vccd1 vccd1 _16533_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13745_ _16297_/Q _13856_/B _13745_/C vssd1 vssd1 vccd1 vccd1 _13745_/Y sky130_fd_sc_hd__nand3_1
X_10957_ _15904_/Q _11183_/B _10963_/C vssd1 vssd1 vccd1 vccd1 _10959_/C sky130_fd_sc_hd__nand3_1
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16464_ input11/X _16464_/D vssd1 vssd1 vccd1 vccd1 _16464_/Q sky130_fd_sc_hd__dfxtp_1
X_13676_ _16289_/Q _13900_/B _13676_/C vssd1 vssd1 vccd1 vccd1 _13676_/X sky130_fd_sc_hd__and3_1
X_10888_ _10888_/A vssd1 vssd1 vccd1 vccd1 _15893_/D sky130_fd_sc_hd__clkbuf_1
X_15415_ _15415_/A vssd1 vssd1 vccd1 vccd1 _15440_/A sky130_fd_sc_hd__clkbuf_4
X_12627_ _16140_/Q _12634_/C _12567_/X vssd1 vssd1 vccd1 vccd1 _12627_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16395_ input11/X _16395_/D vssd1 vssd1 vccd1 vccd1 _16395_/Q sky130_fd_sc_hd__dfxtp_1
X_15346_ _16551_/Q _15346_/B _15346_/C vssd1 vssd1 vccd1 vccd1 _15347_/B sky130_fd_sc_hd__and3_1
X_12558_ _12558_/A vssd1 vssd1 vccd1 vccd1 _16129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ _11737_/A _11509_/B _11509_/C vssd1 vssd1 vccd1 vccd1 _11510_/C sky130_fd_sc_hd__or3_1
X_15277_ _16522_/Q _16521_/Q _16520_/Q _15172_/X vssd1 vssd1 vccd1 vccd1 _16532_/D
+ sky130_fd_sc_hd__o31a_1
X_12489_ _12483_/C _12484_/C _12486_/Y _12487_/X vssd1 vssd1 vccd1 vccd1 _12490_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_144_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14228_ _14342_/A _14228_/B _14232_/A vssd1 vssd1 vccd1 vccd1 _16366_/D sky130_fd_sc_hd__nor3_1
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _14157_/A _14157_/B _14158_/X vssd1 vssd1 vccd1 vccd1 _16356_/D sky130_fd_sc_hd__a21oi_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08720_ _15477_/Q _08721_/C _15335_/B vssd1 vssd1 vccd1 vccd1 _08723_/B sky130_fd_sc_hd__a21o_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08651_ _09038_/A _08705_/B _08651_/C vssd1 vssd1 vccd1 vccd1 _08656_/A sky130_fd_sc_hd__and3_1
XFILLER_82_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08582_ _10956_/A vssd1 vssd1 vccd1 vccd1 _10486_/A sky130_fd_sc_hd__buf_4
XFILLER_93_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09203_ _09203_/A _09203_/B vssd1 vssd1 vccd1 vccd1 _15576_/D sky130_fd_sc_hd__nor2_1
XFILLER_50_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09134_ _09139_/C vssd1 vssd1 vccd1 vccd1 _09150_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_09065_ _15550_/Q _09145_/B _09070_/C vssd1 vssd1 vccd1 vccd1 _09072_/A sky130_fd_sc_hd__and3_1
X_08016_ _14222_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _08222_/B sky130_fd_sc_hd__xnor2_2
XFILLER_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09967_ _15731_/Q _09966_/C _08629_/A vssd1 vssd1 vccd1 vccd1 _09968_/B sky130_fd_sc_hd__a21o_1
XFILLER_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08918_ _09037_/A _08921_/C vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__and2_1
X_09898_ _09898_/A vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__buf_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08849_ _15504_/Q _09016_/B _08849_/C vssd1 vssd1 vccd1 vccd1 _08851_/C sky130_fd_sc_hd__nand3_1
XFILLER_73_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11860_ _16031_/Q _11969_/B _11869_/C vssd1 vssd1 vccd1 vccd1 _11865_/A sky130_fd_sc_hd__and3_1
XFILLER_26_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10811_ _12574_/A vssd1 vssd1 vccd1 vccd1 _10812_/B sky130_fd_sc_hd__buf_2
XFILLER_26_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11791_ _11903_/A vssd1 vssd1 vccd1 vccd1 _11832_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13530_ _16268_/Q _13538_/C _13414_/X vssd1 vssd1 vccd1 vccd1 _13530_/Y sky130_fd_sc_hd__a21oi_1
X_10742_ _15873_/Q _10922_/B _10749_/C vssd1 vssd1 vccd1 vccd1 _10742_/X sky130_fd_sc_hd__and3_1
XFILLER_41_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10673_ _11233_/A vssd1 vssd1 vccd1 vccd1 _10673_/X sky130_fd_sc_hd__buf_2
X_13461_ _13459_/Y _13455_/C _13457_/Y _13458_/X vssd1 vssd1 vccd1 vccd1 _13462_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15200_ _16520_/Q _15209_/C _10797_/B vssd1 vssd1 vccd1 vccd1 _15200_/Y sky130_fd_sc_hd__a21oi_1
X_12412_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12418_/C sky130_fd_sc_hd__nor2_1
XFILLER_138_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16180_ _16555_/Q _16180_/D vssd1 vssd1 vccd1 vccd1 _16180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13392_ _13392_/A vssd1 vssd1 vccd1 vccd1 _13617_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15131_ _15131_/A _15131_/B _15131_/C vssd1 vssd1 vccd1 vccd1 _15132_/C sky130_fd_sc_hd__nand3_1
X_12343_ _12343_/A _12343_/B _12343_/C vssd1 vssd1 vccd1 vccd1 _12344_/A sky130_fd_sc_hd__and3_1
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15062_ _15221_/A vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__clkbuf_2
X_12274_ _12283_/A _12274_/B _12274_/C vssd1 vssd1 vccd1 vccd1 _12275_/A sky130_fd_sc_hd__and3_1
XFILLER_141_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11225_ _13545_/A vssd1 vssd1 vccd1 vccd1 _11452_/A sky130_fd_sc_hd__clkbuf_2
X_14013_ _14035_/A _14013_/B _14013_/C vssd1 vssd1 vccd1 vccd1 _14014_/A sky130_fd_sc_hd__and3_1
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11156_ _11236_/A _11156_/B _11163_/B vssd1 vssd1 vccd1 vccd1 _15931_/D sky130_fd_sc_hd__nor3_1
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10107_ _10107_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10109_/A sky130_fd_sc_hd__or2_1
X_15964_ _16005_/CLK _15964_/D vssd1 vssd1 vccd1 vccd1 _15964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11087_ _11085_/Y _11081_/C _11083_/Y _11084_/X vssd1 vssd1 vccd1 vccd1 _11088_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10038_ _15746_/Q _10190_/B _10038_/C vssd1 vssd1 vccd1 vccd1 _10038_/X sky130_fd_sc_hd__and3_1
X_14915_ _14936_/A _14915_/B _14915_/C vssd1 vssd1 vccd1 vccd1 _14916_/A sky130_fd_sc_hd__and3_1
X_15895_ _16553_/Q _15895_/D vssd1 vssd1 vccd1 vccd1 _15895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14846_ _14881_/C vssd1 vssd1 vccd1 vccd1 _14887_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ _14777_/A vssd1 vssd1 vccd1 vccd1 _15007_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11989_ _11987_/Y _11982_/C _11984_/Y _11986_/X vssd1 vssd1 vccd1 vccd1 _11990_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16516_ _16595_/CLK _16516_/D vssd1 vssd1 vccd1 vccd1 _16516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13728_ input10/X vssd1 vssd1 vccd1 vccd1 _14851_/A sky130_fd_sc_hd__buf_4
XFILLER_32_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16447_ _16607_/CLK _16447_/D vssd1 vssd1 vccd1 vccd1 _16447_/Q sky130_fd_sc_hd__dfxtp_1
X_13659_ _14092_/A vssd1 vssd1 vccd1 vccd1 _13784_/A sky130_fd_sc_hd__buf_2
X_16378_ _16389_/CLK _16378_/D vssd1 vssd1 vccd1 vccd1 _16378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15329_ _15453_/Q _15452_/Q _15451_/Q _15172_/X vssd1 vssd1 vccd1 vccd1 _16543_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ _10393_/A vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__buf_2
XFILLER_59_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09752_ _09749_/X _09747_/B _09751_/Y vssd1 vssd1 vccd1 vccd1 _15685_/D sky130_fd_sc_hd__o21a_1
XFILLER_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08703_ _08644_/X _08705_/C _15312_/A vssd1 vssd1 vccd1 vccd1 _08704_/B sky130_fd_sc_hd__o21ai_1
XFILLER_55_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09683_ _09683_/A vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__buf_2
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16623__28 vssd1 vssd1 vccd1 vccd1 _16623__28/HI _16689_/A sky130_fd_sc_hd__conb_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _08700_/A _08651_/C vssd1 vssd1 vccd1 vccd1 _08634_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08564_/Y _08530_/B _08548_/B _08562_/Y _08555_/Y vssd1 vssd1 vccd1 vccd1
+ _08565_/X sky130_fd_sc_hd__a311o_1
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08496_ _08496_/A _08496_/B vssd1 vssd1 vccd1 vccd1 _08502_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ _09117_/A vssd1 vssd1 vccd1 vccd1 _09117_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ _15561_/Q vssd1 vssd1 vccd1 vccd1 _09057_/C sky130_fd_sc_hd__inv_2
XFILLER_89_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _11097_/A _11010_/B _11014_/A vssd1 vssd1 vccd1 vccd1 _15910_/D sky130_fd_sc_hd__nor3_1
XFILLER_150_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12961_ _12957_/Y _12958_/X _12960_/Y _12955_/C vssd1 vssd1 vccd1 vccd1 _12963_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_46_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14700_ _14707_/A _14700_/B _14700_/C vssd1 vssd1 vccd1 vccd1 _14701_/A sky130_fd_sc_hd__and3_1
X_11912_ _16039_/Q _11950_/C _11802_/X vssd1 vssd1 vccd1 vccd1 _11914_/B sky130_fd_sc_hd__a21oi_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _15791_/CLK _15680_/D vssd1 vssd1 vccd1 vccd1 _15680_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _12907_/A _12892_/B _12892_/C vssd1 vssd1 vccd1 vccd1 _12893_/A sky130_fd_sc_hd__and3_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14631_/A vssd1 vssd1 vccd1 vccd1 _16426_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _16029_/Q _11950_/B _11843_/C vssd1 vssd1 vccd1 vccd1 _11852_/B sky130_fd_sc_hd__and3_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14562_ _14597_/C vssd1 vssd1 vccd1 vccd1 _14603_/C sky130_fd_sc_hd__clkbuf_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11771_/Y _11772_/X _11773_/Y _11767_/C vssd1 vssd1 vccd1 vccd1 _11776_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16346_/CLK _16301_/D vssd1 vssd1 vccd1 vccd1 _16301_/Q sky130_fd_sc_hd__dfxtp_1
X_13513_ _16266_/Q _13623_/B _13514_/C vssd1 vssd1 vccd1 vccd1 _13513_/X sky130_fd_sc_hd__and3_1
X_10725_ _15870_/Q _10755_/C _10673_/X vssd1 vssd1 vccd1 vccd1 _10727_/B sky130_fd_sc_hd__a21oi_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _14777_/A vssd1 vssd1 vccd1 vccd1 _14722_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16232_ _16261_/CLK _16232_/D vssd1 vssd1 vccd1 vccd1 _16232_/Q sky130_fd_sc_hd__dfxtp_1
X_13444_ _16256_/Q _13452_/C _13443_/X vssd1 vssd1 vccd1 vccd1 _13447_/B sky130_fd_sc_hd__a21o_1
X_10656_ _10676_/A _10656_/B _10660_/B vssd1 vssd1 vccd1 vccd1 _15854_/D sky130_fd_sc_hd__nor3_1
XFILLER_139_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16163_ _16237_/CLK _16163_/D vssd1 vssd1 vccd1 vccd1 _16163_/Q sky130_fd_sc_hd__dfxtp_1
X_10587_ _10588_/B _10588_/C _10588_/A vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__a21o_1
X_13375_ _13412_/A _13375_/B _13375_/C vssd1 vssd1 vccd1 vccd1 _13376_/A sky130_fd_sc_hd__and3_1
X_15114_ _15112_/A _15112_/B _15113_/X vssd1 vssd1 vccd1 vccd1 _16503_/D sky130_fd_sc_hd__a21oi_1
X_12326_ _12324_/Y _12325_/X _12320_/C _12321_/C vssd1 vssd1 vccd1 vccd1 _12328_/B
+ sky130_fd_sc_hd__o211ai_1
X_16094_ _16118_/CLK _16094_/D vssd1 vssd1 vccd1 vccd1 _16094_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_108_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15045_ _15045_/A _15045_/B _15045_/C vssd1 vssd1 vccd1 vccd1 _15046_/A sky130_fd_sc_hd__and3_1
XFILLER_114_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12257_ _12257_/A _12257_/B _12257_/C vssd1 vssd1 vccd1 vccd1 _12258_/C sky130_fd_sc_hd__nand3_1
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11208_ _11208_/A _11208_/B _11208_/C vssd1 vssd1 vccd1 vccd1 _11209_/A sky130_fd_sc_hd__and3_1
X_12188_ _12222_/A _12188_/B _12188_/C vssd1 vssd1 vccd1 vccd1 _12189_/A sky130_fd_sc_hd__and3_1
X_11139_ _11137_/Y _11131_/C _11133_/Y _11136_/X vssd1 vssd1 vccd1 vccd1 _11140_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15947_ _15365_/A _15947_/D vssd1 vssd1 vccd1 vccd1 _15947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15878_ _16553_/Q _15878_/D vssd1 vssd1 vccd1 vccd1 _15878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14829_ _16459_/Q _14831_/C _14828_/X vssd1 vssd1 vccd1 vccd1 _14832_/A sky130_fd_sc_hd__a21oi_1
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08350_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08350_/X sky130_fd_sc_hd__and2_1
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08281_ _08094_/A _08094_/B _08280_/Y vssd1 vssd1 vccd1 vccd1 _08400_/B sky130_fd_sc_hd__o21a_1
XFILLER_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09804_ _10900_/B vssd1 vssd1 vccd1 vccd1 _10729_/B sky130_fd_sc_hd__buf_4
X_07996_ _16563_/Q _16561_/Q vssd1 vssd1 vccd1 vccd1 _07997_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09735_ _09734_/X _09733_/Y _09644_/X vssd1 vssd1 vccd1 vccd1 _09735_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09666_ _09669_/C vssd1 vssd1 vccd1 vccd1 _09679_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08617_ _15461_/Q _08619_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _08620_/A sky130_fd_sc_hd__a21oi_1
XFILLER_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09597_ _15658_/Q _09641_/B _09603_/C vssd1 vssd1 vccd1 vccd1 _09599_/B sky130_fd_sc_hd__and3_1
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08555_/A _08548_/B vssd1 vssd1 vccd1 vccd1 _08548_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08479_ _08518_/A _08479_/B vssd1 vssd1 vccd1 vccd1 _08480_/B sky130_fd_sc_hd__or2_1
X_10510_ _10510_/A vssd1 vssd1 vccd1 vccd1 _10702_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11490_ _11488_/Y _11483_/C _11486_/Y _11487_/X vssd1 vssd1 vccd1 vccd1 _11491_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10441_ _10439_/Y _10440_/X _10436_/C _10437_/C vssd1 vssd1 vccd1 vccd1 _10443_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_148_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13160_ _16215_/Q _13383_/B _13171_/C vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__and3_1
X_10372_ _10168_/X _10370_/B _10224_/X vssd1 vssd1 vccd1 vccd1 _10372_/Y sky130_fd_sc_hd__a21oi_1
X_12111_ _12105_/Y _12106_/X _12110_/Y _12103_/C vssd1 vssd1 vccd1 vccd1 _12113_/B
+ sky130_fd_sc_hd__o211ai_1
X_13091_ _13317_/A vssd1 vssd1 vccd1 vccd1 _13131_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12042_ _12042_/A vssd1 vssd1 vccd1 vccd1 _16056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15801_ _15812_/CLK _15801_/D vssd1 vssd1 vccd1 vccd1 _15801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13993_ _14158_/A _13997_/C vssd1 vssd1 vccd1 vccd1 _13993_/X sky130_fd_sc_hd__or2_1
X_15732_ _15812_/CLK _15732_/D vssd1 vssd1 vccd1 vccd1 _15732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _16185_/Q _12952_/C _12887_/X vssd1 vssd1 vccd1 vccd1 _12944_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_65_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15663_ _15791_/CLK _15663_/D vssd1 vssd1 vccd1 vccd1 _15663_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12875_ _16175_/Q _12916_/C _12650_/X vssd1 vssd1 vccd1 vccd1 _12878_/B sky130_fd_sc_hd__a21oi_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14614_ _14614_/A vssd1 vssd1 vccd1 vccd1 _16423_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _16027_/Q _11836_/C _11770_/X vssd1 vssd1 vccd1 vccd1 _11826_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _16551_/CLK _15594_/D vssd1 vssd1 vccd1 vccd1 _15594_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _16414_/Q _14547_/C _14544_/X vssd1 vssd1 vccd1 vccd1 _14548_/A sky130_fd_sc_hd__a21oi_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11757_ _16017_/Q _11922_/B _11757_/C vssd1 vssd1 vccd1 vccd1 _11757_/X sky130_fd_sc_hd__and3_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10708_ _10708_/A _10708_/B vssd1 vssd1 vccd1 vccd1 _10710_/A sky130_fd_sc_hd__or2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14476_ _14476_/A _14476_/B _14476_/C vssd1 vssd1 vccd1 vccd1 _14477_/A sky130_fd_sc_hd__and3_1
X_11688_ _16007_/Q _11688_/B _11698_/C vssd1 vssd1 vccd1 vccd1 _11693_/A sky130_fd_sc_hd__and3_1
X_16215_ _16261_/CLK _16215_/D vssd1 vssd1 vccd1 vccd1 _16215_/Q sky130_fd_sc_hd__dfxtp_1
X_13427_ _13427_/A _13427_/B vssd1 vssd1 vccd1 vccd1 _13432_/C sky130_fd_sc_hd__nor2_1
X_10639_ _15854_/Q _10735_/B _10639_/C vssd1 vssd1 vccd1 vccd1 _10639_/X sky130_fd_sc_hd__and3_1
X_16146_ _16555_/Q _16146_/D vssd1 vssd1 vccd1 vccd1 _16146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _16244_/Q _13586_/B _13358_/C vssd1 vssd1 vccd1 vccd1 _13366_/A sky130_fd_sc_hd__and3_1
XFILLER_142_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ _12332_/C vssd1 vssd1 vccd1 vccd1 _12346_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16077_ _16554_/Q _16077_/D vssd1 vssd1 vccd1 vccd1 _16077_/Q sky130_fd_sc_hd__dfxtp_1
X_13289_ _14411_/A vssd1 vssd1 vccd1 vccd1 _13289_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15028_ _15026_/Y _15027_/X _15023_/C _15024_/C vssd1 vssd1 vccd1 vccd1 _15030_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_69_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07850_ input8/X vssd1 vssd1 vccd1 vccd1 _09278_/A sky130_fd_sc_hd__buf_2
XFILLER_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07781_ input1/X vssd1 vssd1 vccd1 vccd1 _07806_/A sky130_fd_sc_hd__buf_4
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_8
XFILLER_77_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09520_ _15641_/Q _09519_/C _09383_/X vssd1 vssd1 vccd1 vccd1 _09521_/B sky130_fd_sc_hd__a21o_1
XFILLER_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09451_ _15629_/Q _09585_/B _09458_/C vssd1 vssd1 vccd1 vccd1 _09453_/C sky130_fd_sc_hd__nand3_1
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08402_ _08469_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08403_/B sky130_fd_sc_hd__xor2_4
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09382_ _15614_/Q _09472_/B _09382_/C vssd1 vssd1 vccd1 vccd1 _09382_/X sky130_fd_sc_hd__and3_1
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08333_ _08333_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08333_/Y sky130_fd_sc_hd__nor2_1
X_08264_ _08590_/C _15335_/C _08263_/Y vssd1 vssd1 vccd1 vccd1 _08385_/C sky130_fd_sc_hd__o21ai_4
X_08195_ _08195_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08323_/A sky130_fd_sc_hd__xnor2_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _16577_/Q vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__inv_2
XFILLER_142_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09718_ _09718_/A _09718_/B _09722_/A vssd1 vssd1 vccd1 vccd1 _15679_/D sky130_fd_sc_hd__nor3_1
XFILLER_74_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10990_ _11097_/A _10990_/B _10994_/B vssd1 vssd1 vccd1 vccd1 _15907_/D sky130_fd_sc_hd__nor3_1
XFILLER_43_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09649_ _15668_/Q _09648_/C _09604_/X vssd1 vssd1 vccd1 vccd1 _09650_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12681_/A _12660_/B _12660_/C vssd1 vssd1 vccd1 vccd1 _12661_/A sky130_fd_sc_hd__and3_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11666_/A _11611_/B _11615_/B vssd1 vssd1 vccd1 vccd1 _15995_/D sky130_fd_sc_hd__nor3_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12591_ _12614_/C vssd1 vssd1 vccd1 vccd1 _12628_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ _14332_/B _14332_/C _14108_/X vssd1 vssd1 vccd1 vccd1 _14333_/B sky130_fd_sc_hd__o21ai_1
XFILLER_129_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _15987_/Q _11654_/B _11551_/C vssd1 vssd1 vccd1 vccd1 _11542_/X sky130_fd_sc_hd__and3_1
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14261_ _16371_/Q _14318_/B _14268_/C vssd1 vssd1 vccd1 vccd1 _14261_/Y sky130_fd_sc_hd__nand3_1
X_11473_ _15977_/Q _11638_/B _11473_/C vssd1 vssd1 vccd1 vccd1 _11473_/X sky130_fd_sc_hd__and3_1
X_16000_ _16005_/CLK _16000_/D vssd1 vssd1 vccd1 vccd1 _16000_/Q sky130_fd_sc_hd__dfxtp_1
X_13212_ _13212_/A vssd1 vssd1 vccd1 vccd1 _13228_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10424_ _10440_/C vssd1 vssd1 vccd1 vccd1 _10457_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14192_ _16363_/Q _14201_/C _14029_/X vssd1 vssd1 vccd1 vccd1 _14192_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_136_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13143_ _16213_/Q _13364_/B _13143_/C vssd1 vssd1 vccd1 vccd1 _13151_/B sky130_fd_sc_hd__and3_1
XFILLER_136_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10355_ _15802_/Q _10402_/B _10355_/C vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__and3_1
XFILLER_3_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16659__64 vssd1 vssd1 vccd1 vccd1 _16659__64/HI _16735_/A sky130_fd_sc_hd__conb_1
X_10286_ _10311_/A _10286_/B _10290_/A vssd1 vssd1 vccd1 vccd1 _15787_/D sky130_fd_sc_hd__nor3_1
X_13074_ _16204_/Q _13082_/C _12850_/X vssd1 vssd1 vccd1 vccd1 _13074_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12025_ _16055_/Q _12065_/C _11802_/X vssd1 vssd1 vccd1 vccd1 _12028_/B sky130_fd_sc_hd__a21oi_1
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13976_ _13974_/Y _13969_/C _13971_/Y _13973_/X vssd1 vssd1 vccd1 vccd1 _13977_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_46_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15715_ _15812_/CLK _15715_/D vssd1 vssd1 vccd1 vccd1 _15715_/Q sky130_fd_sc_hd__dfxtp_2
X_12927_ _12927_/A vssd1 vssd1 vccd1 vccd1 _16181_/D sky130_fd_sc_hd__clkbuf_1
X_16695_ _16695_/A _07793_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_34_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15646_ _15791_/CLK _15646_/D vssd1 vssd1 vccd1 vccd1 _15646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12858_ _16173_/Q _12860_/C _12857_/X vssd1 vssd1 vccd1 vccd1 _12861_/A sky130_fd_sc_hd__a21oi_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ _11810_/B _11810_/C _11810_/A vssd1 vssd1 vccd1 vccd1 _11811_/B sky130_fd_sc_hd__a21o_1
X_15577_ _16551_/CLK _15577_/D vssd1 vssd1 vccd1 vccd1 _15577_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12789_/A vssd1 vssd1 vccd1 vccd1 _16162_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14528_ _14528_/A vssd1 vssd1 vccd1 vccd1 _16410_/D sky130_fd_sc_hd__clkbuf_1
X_14459_ _14457_/Y _14458_/X _14454_/C _14455_/C vssd1 vssd1 vccd1 vccd1 _14461_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_128_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16129_ _16554_/Q _16129_/D vssd1 vssd1 vccd1 vccd1 _16129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08951_ _08951_/A _08951_/B vssd1 vssd1 vccd1 vccd1 _08952_/B sky130_fd_sc_hd__nor2_1
XFILLER_142_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07902_ _15678_/Q vssd1 vssd1 vccd1 vccd1 _09625_/C sky130_fd_sc_hd__clkinv_4
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08882_ _08882_/A _08882_/B vssd1 vssd1 vccd1 vccd1 _15505_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07833_ _07836_/A vssd1 vssd1 vccd1 vccd1 _07833_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07764_ _07768_/A vssd1 vssd1 vccd1 vccd1 _07764_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09503_ _09503_/A vssd1 vssd1 vccd1 vccd1 _15635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09434_ _09427_/Y _09428_/X _09430_/B vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__o21a_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09365_ _09366_/B _09366_/C _09366_/A vssd1 vssd1 vccd1 vccd1 _09367_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08316_ _08316_/A _08301_/A vssd1 vssd1 vccd1 vccd1 _08413_/A sky130_fd_sc_hd__or2b_1
X_09296_ _09436_/A _09296_/B vssd1 vssd1 vccd1 vccd1 _09296_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_30 _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ _15013_/A _08247_/B vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__or2_1
XFILLER_20_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08178_ _16578_/Q _08178_/B vssd1 vssd1 vccd1 vccd1 _08178_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10140_ _15765_/Q _10300_/C _10152_/C vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__and3_1
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10071_ _10578_/A vssd1 vssd1 vccd1 vccd1 _10179_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13830_ _13831_/B _13831_/C _13829_/X vssd1 vssd1 vccd1 vccd1 _13832_/B sky130_fd_sc_hd__o21ai_1
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ _13758_/Y _13767_/A _13760_/Y _13756_/C vssd1 vssd1 vccd1 vccd1 _13763_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10973_ _10981_/A _10973_/B _10973_/C vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__and3_1
X_15500_ _16551_/CLK _15500_/D vssd1 vssd1 vccd1 vccd1 _15500_/Q sky130_fd_sc_hd__dfxtp_2
X_12712_ _16152_/Q _12881_/B _12718_/C vssd1 vssd1 vccd1 vccd1 _12714_/C sky130_fd_sc_hd__nand3_1
XFILLER_16_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _16607_/CLK _16480_/D vssd1 vssd1 vccd1 vccd1 _16480_/Q sky130_fd_sc_hd__dfxtp_1
X_13692_ _16291_/Q _13914_/B _13700_/C vssd1 vssd1 vccd1 vccd1 _13692_/X sky130_fd_sc_hd__and3_1
X_15431_ _16293_/Q _16292_/Q _16291_/Q _15428_/X vssd1 vssd1 vccd1 vccd1 _16607_/D
+ sky130_fd_sc_hd__o31a_1
X_12643_ _12868_/A _12643_/B _12643_/C vssd1 vssd1 vccd1 vccd1 _12644_/C sky130_fd_sc_hd__or3_1
XFILLER_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15362_ _08663_/X _15360_/A _15361_/Y vssd1 vssd1 vccd1 vccd1 _16551_/D sky130_fd_sc_hd__o21a_1
X_12574_ _12574_/A vssd1 vssd1 vccd1 vccd1 _13705_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14313_ _14311_/Y _14306_/C _14309_/Y _14310_/X vssd1 vssd1 vccd1 vccd1 _14314_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11525_ _11525_/A _11525_/B _11525_/C vssd1 vssd1 vccd1 vccd1 _11526_/C sky130_fd_sc_hd__nand3_1
X_15293_ _16706_/A _15306_/A _15293_/C vssd1 vssd1 vccd1 vccd1 _15293_/X sky130_fd_sc_hd__and3_1
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14244_ _16370_/Q _14464_/B _14245_/C vssd1 vssd1 vccd1 vccd1 _14244_/X sky130_fd_sc_hd__and3_1
X_11456_ _11473_/C vssd1 vssd1 vccd1 vccd1 _11480_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10407_ _15812_/Q _10408_/C _10360_/X vssd1 vssd1 vccd1 vccd1 _10409_/A sky130_fd_sc_hd__a21oi_1
X_14175_ _14175_/A _14175_/B _14175_/C vssd1 vssd1 vccd1 vccd1 _14176_/C sky130_fd_sc_hd__nand3_1
X_11387_ _11385_/A _11385_/B _11386_/X vssd1 vssd1 vccd1 vccd1 _15964_/D sky130_fd_sc_hd__a21oi_1
XFILLER_125_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13126_ _13407_/A vssd1 vssd1 vccd1 vccd1 _13350_/B sky130_fd_sc_hd__clkbuf_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ _10338_/A _10338_/B _10338_/C vssd1 vssd1 vccd1 vccd1 _10339_/A sky130_fd_sc_hd__and3_1
XFILLER_98_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13057_/A vssd1 vssd1 vccd1 vccd1 _16200_/D sky130_fd_sc_hd__clkbuf_1
X_10269_ _10269_/A _10269_/B vssd1 vssd1 vccd1 vccd1 _10270_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ _16053_/Q _12010_/C _12007_/X vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__a21oi_1
XFILLER_94_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13959_ _13956_/Y _13958_/X _13953_/C _13954_/C vssd1 vssd1 vccd1 vccd1 _13961_/B
+ sky130_fd_sc_hd__o211ai_1
X_16747_ _16747_/A _07764_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15629_ _15791_/CLK _15629_/D vssd1 vssd1 vccd1 vccd1 _15629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09150_ _15569_/Q _09192_/B _09150_/C vssd1 vssd1 vccd1 vccd1 _09151_/B sky130_fd_sc_hd__and3_1
X_08101_ _15534_/Q _08114_/B vssd1 vssd1 vccd1 vccd1 _08102_/B sky130_fd_sc_hd__xnor2_2
XFILLER_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09081_ _09240_/A _09084_/C vssd1 vssd1 vccd1 vccd1 _09083_/A sky130_fd_sc_hd__and2_1
XFILLER_147_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08032_ _15795_/Q _15777_/Q vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ _15722_/Q _15721_/Q _15720_/Q _09982_/X vssd1 vssd1 vccd1 vccd1 _15732_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_103_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08934_ _15521_/Q _09053_/B _08937_/C vssd1 vssd1 vccd1 vccd1 _08939_/A sky130_fd_sc_hd__and3_1
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08865_ _15506_/Q _08866_/C _08777_/X vssd1 vssd1 vccd1 vccd1 _08867_/A sky130_fd_sc_hd__a21oi_1
XFILLER_85_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07816_ _07818_/A vssd1 vssd1 vccd1 vccd1 _07816_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08796_ _09207_/A vssd1 vssd1 vccd1 vccd1 _08796_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09417_ _09415_/Y _09422_/A _09412_/C _09413_/C vssd1 vssd1 vccd1 vccd1 _09419_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09348_ _09291_/X _09346_/B _09347_/Y vssd1 vssd1 vccd1 vccd1 _15603_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09279_ _09698_/A vssd1 vssd1 vccd1 vccd1 _10017_/A sky130_fd_sc_hd__buf_2
XFILLER_148_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _11307_/Y _11308_/X _11309_/Y _11304_/C vssd1 vssd1 vccd1 vccd1 _11312_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_126_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12290_ _12288_/Y _12283_/C _12286_/Y _12298_/A vssd1 vssd1 vccd1 vccd1 _12298_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11241_ _11242_/B _11242_/C _11242_/A vssd1 vssd1 vccd1 vccd1 _11243_/B sky130_fd_sc_hd__a21o_1
XFILLER_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11172_ _16563_/Q vssd1 vssd1 vccd1 vccd1 _11190_/C sky130_fd_sc_hd__inv_2
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _15762_/Q _10158_/C _09943_/X vssd1 vssd1 vccd1 vccd1 _10125_/B sky130_fd_sc_hd__a21oi_1
X_16629__34 vssd1 vssd1 vccd1 vccd1 _16629__34/HI _16695_/A sky130_fd_sc_hd__conb_1
X_15980_ _16005_/CLK _15980_/D vssd1 vssd1 vccd1 vccd1 _15980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10054_ _10052_/Y _10048_/C _10050_/Y _10059_/A vssd1 vssd1 vccd1 vccd1 _10059_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14931_ _16475_/Q _15041_/B _14940_/C vssd1 vssd1 vccd1 vccd1 _14931_/X sky130_fd_sc_hd__and3_1
XFILLER_57_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14862_ _14855_/C _14856_/C _14859_/Y _14860_/X vssd1 vssd1 vccd1 vccd1 _14863_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16601_ _16607_/CLK _16601_/D vssd1 vssd1 vccd1 vccd1 _16601_/Q sky130_fd_sc_hd__dfxtp_1
X_13813_ _14092_/A vssd1 vssd1 vccd1 vccd1 _13927_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14793_ _16454_/Q _14853_/B _14800_/C vssd1 vssd1 vccd1 vccd1 _14795_/C sky130_fd_sc_hd__nand3_1
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16532_ _16595_/CLK _16532_/D vssd1 vssd1 vccd1 vccd1 _16532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13744_ _16298_/Q _13906_/B _13745_/C vssd1 vssd1 vccd1 vccd1 _13744_/X sky130_fd_sc_hd__and3_1
X_10956_ _10956_/A vssd1 vssd1 vccd1 vccd1 _11183_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_44_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16463_ input11/X _16463_/D vssd1 vssd1 vccd1 vccd1 _16463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13675_ _14799_/A vssd1 vssd1 vccd1 vccd1 _13900_/B sky130_fd_sc_hd__clkbuf_2
X_10887_ _10925_/A _10887_/B _10887_/C vssd1 vssd1 vccd1 vccd1 _10888_/A sky130_fd_sc_hd__and3_1
X_15414_ _16189_/Q _16188_/Q _16187_/Q _15409_/X vssd1 vssd1 vccd1 vccd1 _16594_/D
+ sky130_fd_sc_hd__o31a_1
X_12626_ _12626_/A vssd1 vssd1 vccd1 vccd1 _16138_/D sky130_fd_sc_hd__clkbuf_1
X_16394_ input11/X _16394_/D vssd1 vssd1 vccd1 vccd1 _16394_/Q sky130_fd_sc_hd__dfxtp_1
X_15345_ _16551_/Q _15346_/C _10510_/A vssd1 vssd1 vccd1 vccd1 _15347_/A sky130_fd_sc_hd__a21oi_1
X_12557_ _12565_/A _12557_/B _12557_/C vssd1 vssd1 vccd1 vccd1 _12558_/A sky130_fd_sc_hd__and3_1
XFILLER_129_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11508_ _13545_/A vssd1 vssd1 vccd1 vccd1 _11737_/A sky130_fd_sc_hd__clkbuf_2
X_15276_ _15276_/A vssd1 vssd1 vccd1 vccd1 _16531_/D sky130_fd_sc_hd__clkbuf_1
X_12488_ _12486_/Y _12487_/X _12483_/C _12484_/C vssd1 vssd1 vccd1 vccd1 _12490_/B
+ sky130_fd_sc_hd__o211ai_1
X_14227_ _16367_/Q _14227_/B _14237_/C vssd1 vssd1 vccd1 vccd1 _14232_/A sky130_fd_sc_hd__and3_1
X_11439_ _11437_/Y _11431_/C _11435_/Y _11446_/A vssd1 vssd1 vccd1 vccd1 _11446_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_113_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14158_ _14158_/A _14162_/C vssd1 vssd1 vccd1 vccd1 _14158_/X sky130_fd_sc_hd__or2_1
XFILLER_113_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _13109_/A vssd1 vssd1 vccd1 vccd1 _16207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _14087_/Y _14082_/C _14084_/Y _14085_/X vssd1 vssd1 vccd1 vccd1 _14090_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_79_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08650_ _09164_/A vssd1 vssd1 vccd1 vccd1 _08705_/B sky130_fd_sc_hd__buf_2
XFILLER_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08581_ _12655_/A vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__buf_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _09038_/X _09204_/C _09126_/X vssd1 vssd1 vccd1 vccd1 _09203_/B sky130_fd_sc_hd__o21ai_1
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ _15579_/Q vssd1 vssd1 vccd1 vccd1 _09139_/C sky130_fd_sc_hd__inv_2
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09064_ _15550_/Q _09070_/C _09063_/X vssd1 vssd1 vccd1 vccd1 _09064_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08015_ _14335_/A _08214_/B vssd1 vssd1 vccd1 vccd1 _08016_/B sky130_fd_sc_hd__xnor2_2
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09966_ _15731_/Q _09966_/B _09966_/C vssd1 vssd1 vccd1 vccd1 _09966_/X sky130_fd_sc_hd__and3_1
XFILLER_134_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08917_ _08872_/X _08908_/B _08912_/B _08916_/Y vssd1 vssd1 vccd1 vccd1 _15512_/D
+ sky130_fd_sc_hd__o31a_1
X_09897_ _08654_/X _09891_/B _09792_/X vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__a21oi_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08848_ _09056_/A vssd1 vssd1 vccd1 vccd1 _09016_/B sky130_fd_sc_hd__buf_2
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08779_ _15488_/Q _09271_/A _08779_/C vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__and3_1
X_10810_ _15884_/Q _10812_/C _09164_/A vssd1 vssd1 vccd1 vccd1 _10813_/A sky130_fd_sc_hd__a21oi_1
XFILLER_25_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11790_ _11788_/A _11788_/B _11789_/X vssd1 vssd1 vccd1 vccd1 _16020_/D sky130_fd_sc_hd__a21oi_1
X_10741_ _15873_/Q _10749_/C _09683_/A vssd1 vssd1 vccd1 vccd1 _10741_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ _13457_/Y _13458_/X _13459_/Y _13455_/C vssd1 vssd1 vccd1 vccd1 _13462_/B
+ sky130_fd_sc_hd__o211ai_1
X_10672_ _10701_/C vssd1 vssd1 vccd1 vccd1 _10707_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12411_ _12411_/A _12411_/B vssd1 vssd1 vccd1 vccd1 _12412_/B sky130_fd_sc_hd__nor2_1
X_13391_ _16249_/Q _13401_/C _13169_/X vssd1 vssd1 vccd1 vccd1 _13391_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15130_ _15131_/B _15131_/C _15131_/A vssd1 vssd1 vccd1 vccd1 _15132_/B sky130_fd_sc_hd__a21o_1
XFILLER_127_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12342_ _12340_/Y _12335_/C _12338_/Y _12339_/X vssd1 vssd1 vccd1 vccd1 _12343_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15061_ _15059_/A _15059_/B _15060_/X vssd1 vssd1 vccd1 vccd1 _16494_/D sky130_fd_sc_hd__a21oi_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ _12271_/Y _12266_/C _12268_/Y _12270_/X vssd1 vssd1 vccd1 vccd1 _12274_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14012_ _14012_/A _14012_/B _14012_/C vssd1 vssd1 vccd1 vccd1 _14013_/C sky130_fd_sc_hd__nand3_1
X_11224_ _11226_/B _11226_/C _10999_/X vssd1 vssd1 vccd1 vccd1 _11227_/B sky130_fd_sc_hd__o21ai_1
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11155_ _11153_/Y _11148_/C _11151_/Y _11163_/A vssd1 vssd1 vccd1 vccd1 _11163_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_49_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10106_ _15758_/Q _10313_/C _10106_/C vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__and3_1
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15963_ _16005_/CLK _15963_/D vssd1 vssd1 vccd1 vccd1 _15963_/Q sky130_fd_sc_hd__dfxtp_1
X_11086_ _11083_/Y _11084_/X _11085_/Y _11081_/C vssd1 vssd1 vccd1 vccd1 _11088_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_76_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10037_ _15746_/Q _10038_/C _09813_/X vssd1 vssd1 vccd1 vccd1 _10037_/Y sky130_fd_sc_hd__a21oi_1
X_14914_ _14914_/A _14914_/B _14914_/C vssd1 vssd1 vccd1 vccd1 _14915_/C sky130_fd_sc_hd__nand3_1
XFILLER_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15894_ _16553_/Q _15894_/D vssd1 vssd1 vccd1 vccd1 _15894_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14845_ _14867_/C vssd1 vssd1 vccd1 vccd1 _14881_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14776_ _14774_/A _14774_/B _14775_/X vssd1 vssd1 vccd1 vccd1 _16449_/D sky130_fd_sc_hd__a21oi_1
X_11988_ _11984_/Y _11986_/X _11987_/Y _11982_/C vssd1 vssd1 vccd1 vccd1 _11990_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13727_ _13784_/A _13727_/B _13733_/A vssd1 vssd1 vccd1 vccd1 _16294_/D sky130_fd_sc_hd__nor3_1
X_16515_ _16607_/CLK _16515_/D vssd1 vssd1 vccd1 vccd1 _16515_/Q sky130_fd_sc_hd__dfxtp_2
X_10939_ _10937_/A _10937_/B _10938_/X vssd1 vssd1 vccd1 vccd1 _15900_/D sky130_fd_sc_hd__a21oi_1
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16446_ _16607_/CLK _16446_/D vssd1 vssd1 vccd1 vccd1 _16446_/Q sky130_fd_sc_hd__dfxtp_1
X_13658_ _13658_/A vssd1 vssd1 vccd1 vccd1 _16285_/D sky130_fd_sc_hd__clkbuf_1
X_12609_ _12602_/C _12603_/C _12606_/Y _12607_/X vssd1 vssd1 vccd1 vccd1 _12610_/C
+ sky130_fd_sc_hd__a211o_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16377_ _16389_/CLK _16377_/D vssd1 vssd1 vccd1 vccd1 _16377_/Q sky130_fd_sc_hd__dfxtp_1
X_13589_ _13587_/Y _13583_/C _13585_/Y _13594_/A vssd1 vssd1 vccd1 vccd1 _13594_/B
+ sky130_fd_sc_hd__a211oi_1
X_15328_ _08567_/X _15327_/X _15325_/X _15367_/B vssd1 vssd1 vccd1 vccd1 _16542_/D
+ sky130_fd_sc_hd__a31oi_1
XFILLER_144_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15259_ _15259_/A vssd1 vssd1 vccd1 vccd1 _16528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09820_ _09820_/A vssd1 vssd1 vccd1 vccd1 _15699_/D sky130_fd_sc_hd__clkbuf_1
X_09751_ _09658_/X _09747_/B _09750_/X vssd1 vssd1 vccd1 vccd1 _09751_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08702_ _08831_/A _08705_/C vssd1 vssd1 vccd1 vccd1 _08704_/A sky130_fd_sc_hd__and2_1
X_09682_ _09718_/A _09682_/B _09687_/B vssd1 vssd1 vccd1 vccd1 _15672_/D sky130_fd_sc_hd__nor3_1
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08633_ _08620_/B _08623_/B _09076_/A vssd1 vssd1 vccd1 vccd1 _08651_/C sky130_fd_sc_hd__o21a_1
XFILLER_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _08564_/A vssd1 vssd1 vccd1 vccd1 _08564_/Y sky130_fd_sc_hd__inv_2
X_08495_ _08445_/A _08445_/B _08494_/X vssd1 vssd1 vccd1 vccd1 _08515_/A sky130_fd_sc_hd__a21bo_2
XFILLER_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09116_ _09114_/A _09114_/B _09115_/X vssd1 vssd1 vccd1 vccd1 _15556_/D sky130_fd_sc_hd__a21oi_1
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09047_ _15533_/Q _15532_/Q _15531_/Q _08887_/X vssd1 vssd1 vccd1 vccd1 _15543_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ _09950_/B _09950_/C _09950_/A vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__a21o_1
XFILLER_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12960_ _16186_/Q _13187_/B _12967_/C vssd1 vssd1 vccd1 vccd1 _12960_/Y sky130_fd_sc_hd__nand3_1
XFILLER_85_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11911_ _11944_/C vssd1 vssd1 vccd1 vccd1 _11950_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_73_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12891_ _12883_/C _12884_/C _12888_/Y _12889_/X vssd1 vssd1 vccd1 vccd1 _12892_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14651_/A _14630_/B _14630_/C vssd1 vssd1 vccd1 vccd1 _14631_/A sky130_fd_sc_hd__and3_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _16029_/Q _11843_/C _11726_/X vssd1 vssd1 vccd1 vccd1 _11844_/A sky130_fd_sc_hd__a21oi_1
XFILLER_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14583_/C vssd1 vssd1 vccd1 vccd1 _14597_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _16018_/Q _11773_/B _11779_/C vssd1 vssd1 vccd1 vccd1 _11773_/Y sky130_fd_sc_hd__nand3_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16346_/CLK _16300_/D vssd1 vssd1 vccd1 vccd1 _16300_/Q sky130_fd_sc_hd__dfxtp_1
X_13512_ _16266_/Q _13514_/C _13289_/X vssd1 vssd1 vccd1 vccd1 _13512_/Y sky130_fd_sc_hd__a21oi_1
X_10724_ _10749_/C vssd1 vssd1 vccd1 vccd1 _10755_/C sky130_fd_sc_hd__clkbuf_2
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14490_/A _14490_/B _14491_/X vssd1 vssd1 vccd1 vccd1 _16404_/D sky130_fd_sc_hd__a21oi_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _16261_/CLK _16231_/D vssd1 vssd1 vccd1 vccd1 _16231_/Q sky130_fd_sc_hd__dfxtp_1
X_13443_ _13443_/A vssd1 vssd1 vccd1 vccd1 _13443_/X sky130_fd_sc_hd__clkbuf_2
X_10655_ _10653_/Y _10649_/C _10651_/Y _10660_/A vssd1 vssd1 vccd1 vccd1 _10660_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16162_ _16237_/CLK _16162_/D vssd1 vssd1 vccd1 vccd1 _16162_/Q sky130_fd_sc_hd__dfxtp_1
X_13374_ _13432_/A _13374_/B _13374_/C vssd1 vssd1 vccd1 vccd1 _13375_/C sky130_fd_sc_hd__or3_1
XFILLER_139_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10586_ _15844_/Q _10679_/B _10593_/C vssd1 vssd1 vccd1 vccd1 _10588_/C sky130_fd_sc_hd__nand3_1
XFILLER_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15113_ _15271_/A _15117_/C vssd1 vssd1 vccd1 vccd1 _15113_/X sky130_fd_sc_hd__or2_1
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12325_ _16097_/Q _12487_/B _12325_/C vssd1 vssd1 vccd1 vccd1 _12325_/X sky130_fd_sc_hd__and3_1
X_16093_ _16554_/Q _16093_/D vssd1 vssd1 vccd1 vccd1 _16093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15044_ _15042_/Y _15038_/C _15040_/Y _15041_/X vssd1 vssd1 vccd1 vccd1 _15045_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_5_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12256_ _12257_/B _12257_/C _12257_/A vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__a21o_1
XFILLER_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11207_ _11205_/Y _11200_/C _11203_/Y _11204_/X vssd1 vssd1 vccd1 vccd1 _11208_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_123_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12187_ _12304_/A _12187_/B _12187_/C vssd1 vssd1 vccd1 vccd1 _12188_/C sky130_fd_sc_hd__or3_1
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11138_ _11133_/Y _11136_/X _11137_/Y _11131_/C vssd1 vssd1 vccd1 vccd1 _11140_/B
+ sky130_fd_sc_hd__o211ai_1
X_15946_ _15365_/A _15946_/D vssd1 vssd1 vccd1 vccd1 _15946_/Q sky130_fd_sc_hd__dfxtp_1
X_11069_ _15921_/Q _11078_/C _10905_/X vssd1 vssd1 vccd1 vccd1 _11069_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15877_ _16553_/Q _15877_/D vssd1 vssd1 vccd1 vccd1 _15877_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14828_ _14828_/A vssd1 vssd1 vccd1 vccd1 _14828_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14759_ _14757_/Y _14753_/C _14755_/Y _14756_/X vssd1 vssd1 vccd1 vccd1 _14760_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08280_ _15804_/Q _08280_/B vssd1 vssd1 vccd1 vccd1 _08280_/Y sky130_fd_sc_hd__nand2_1
X_16429_ _16595_/CLK _16429_/D vssd1 vssd1 vccd1 vccd1 _16429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09803_ _09841_/A _09803_/B _09809_/A vssd1 vssd1 vccd1 vccd1 _15697_/D sky130_fd_sc_hd__nor3_1
XFILLER_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07995_ _16563_/Q _16561_/Q vssd1 vssd1 vccd1 vccd1 _07997_/A sky130_fd_sc_hd__or2_1
XFILLER_87_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09734_ _09734_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09734_/X sky130_fd_sc_hd__or2_1
XFILLER_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ _15687_/Q vssd1 vssd1 vccd1 vccd1 _09669_/C sky130_fd_sc_hd__inv_2
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ _15346_/B vssd1 vssd1 vccd1 vccd1 _08616_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09596_ _15658_/Q _09603_/C _09463_/X vssd1 vssd1 vccd1 vccd1 _09599_/A sky130_fd_sc_hd__a21oi_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _15452_/Q _08561_/B _15315_/C vssd1 vssd1 vccd1 vccd1 _08548_/B sky130_fd_sc_hd__nand3_1
XFILLER_24_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08478_ _08518_/A _08479_/B vssd1 vssd1 vccd1 vccd1 _08480_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10440_ _15818_/Q _10494_/B _10440_/C vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__and3_1
XFILLER_136_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _10220_/X _10363_/B _10366_/B _10370_/Y vssd1 vssd1 vccd1 vccd1 _15802_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_124_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12110_ _16066_/Q _12340_/B _12118_/C vssd1 vssd1 vccd1 vccd1 _12110_/Y sky130_fd_sc_hd__nand3_1
XFILLER_136_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13090_ _13371_/A vssd1 vssd1 vccd1 vccd1 _13317_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12041_ _12056_/A _12041_/B _12041_/C vssd1 vssd1 vccd1 vccd1 _12042_/A sky130_fd_sc_hd__and3_1
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15800_ _15812_/CLK _15800_/D vssd1 vssd1 vccd1 vccd1 _15800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13992_ _13992_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13997_/C sky130_fd_sc_hd__nor2_1
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15731_ _15812_/CLK _15731_/D vssd1 vssd1 vccd1 vccd1 _15731_/Q sky130_fd_sc_hd__dfxtp_1
X_12943_ _12943_/A vssd1 vssd1 vccd1 vccd1 _16183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15662_ _15791_/CLK _15662_/D vssd1 vssd1 vccd1 vccd1 _15662_/Q sky130_fd_sc_hd__dfxtp_2
X_12874_ _12910_/C vssd1 vssd1 vccd1 vccd1 _12916_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _11825_/A vssd1 vssd1 vccd1 vccd1 _16025_/D sky130_fd_sc_hd__clkbuf_1
X_14613_ _14651_/A _14613_/B _14613_/C vssd1 vssd1 vccd1 vccd1 _14614_/A sky130_fd_sc_hd__and3_1
X_15593_ _16570_/CLK _15593_/D vssd1 vssd1 vccd1 vccd1 _15593_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14544_ _14828_/A vssd1 vssd1 vccd1 vccd1 _14544_/X sky130_fd_sc_hd__buf_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _16017_/Q _11764_/C _11755_/X vssd1 vssd1 vccd1 vccd1 _11756_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10707_ _15866_/Q _10707_/B _10707_/C vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__and3_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14475_ _14473_/Y _14469_/C _14471_/Y _14472_/X vssd1 vssd1 vccd1 vccd1 _14476_/C
+ sky130_fd_sc_hd__a211o_1
X_11687_ _16007_/Q _11729_/C _11517_/X vssd1 vssd1 vccd1 vccd1 _11689_/B sky130_fd_sc_hd__a21oi_1
X_16214_ _16261_/CLK _16214_/D vssd1 vssd1 vccd1 vccd1 _16214_/Q sky130_fd_sc_hd__dfxtp_2
X_13426_ _13426_/A _13426_/B vssd1 vssd1 vccd1 vccd1 _13427_/B sky130_fd_sc_hd__nor2_1
X_10638_ _15854_/Q _10639_/C _10492_/X vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16145_ _16555_/Q _16145_/D vssd1 vssd1 vccd1 vccd1 _16145_/Q sky130_fd_sc_hd__dfxtp_1
X_13357_ _13638_/A vssd1 vssd1 vccd1 vccd1 _13586_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10569_ _10569_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10570_/B sky130_fd_sc_hd__nor2_1
XFILLER_127_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ _12325_/C vssd1 vssd1 vccd1 vccd1 _12332_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16076_ _16554_/Q _16076_/D vssd1 vssd1 vccd1 vccd1 _16076_/Q sky130_fd_sc_hd__dfxtp_1
X_13288_ _13288_/A vssd1 vssd1 vccd1 vccd1 _14411_/A sky130_fd_sc_hd__buf_6
XFILLER_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15027_ _16491_/Q _15027_/B _15027_/C vssd1 vssd1 vccd1 vccd1 _15027_/X sky130_fd_sc_hd__and3_1
XFILLER_142_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12239_ _13652_/A vssd1 vssd1 vccd1 vccd1 _13371_/A sky130_fd_sc_hd__buf_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07780_ _07780_/A vssd1 vssd1 vccd1 vccd1 _07780_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
X_15929_ _16005_/CLK _15929_/D vssd1 vssd1 vccd1 vccd1 _15929_/Q sky130_fd_sc_hd__dfxtp_1
X_09450_ _15629_/Q _09458_/C _09362_/X vssd1 vssd1 vccd1 vccd1 _09453_/B sky130_fd_sc_hd__a21o_1
XFILLER_92_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08401_ _08283_/A _08283_/B _08400_/Y vssd1 vssd1 vccd1 vccd1 _08469_/B sky130_fd_sc_hd__a21oi_2
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09381_ _09378_/A _09377_/Y _09378_/B vssd1 vssd1 vccd1 vccd1 _09381_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08332_ _08332_/A vssd1 vssd1 vccd1 vccd1 _08333_/A sky130_fd_sc_hd__inv_2
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08263_ _15489_/Q _08263_/B vssd1 vssd1 vccd1 vccd1 _08263_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08194_ _08194_/A _08194_/B vssd1 vssd1 vccd1 vccd1 _08195_/B sky130_fd_sc_hd__xor2_4
XFILLER_146_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ _16613_/Q vssd1 vssd1 vccd1 vccd1 _14000_/A sky130_fd_sc_hd__inv_4
XFILLER_28_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09717_ _15682_/Q _09945_/B _09717_/C vssd1 vssd1 vccd1 vccd1 _09722_/A sky130_fd_sc_hd__and3_1
XFILLER_19_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ _15668_/Q _09692_/B _09648_/C vssd1 vssd1 vccd1 vccd1 _09648_/X sky130_fd_sc_hd__and3_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09592_/C vssd1 vssd1 vccd1 vccd1 _09603_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11608_/Y _11604_/C _11606_/Y _11615_/A vssd1 vssd1 vccd1 vccd1 _11615_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12607_/C vssd1 vssd1 vccd1 vccd1 _12614_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11541_ _15987_/Q _11551_/C _11485_/X vssd1 vssd1 vccd1 vccd1 _11541_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ _16372_/Q _14427_/B _14260_/C vssd1 vssd1 vccd1 vccd1 _14270_/A sky130_fd_sc_hd__and3_1
X_11472_ _15977_/Q _11480_/C _11471_/X vssd1 vssd1 vccd1 vccd1 _11472_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13211_ _13211_/A vssd1 vssd1 vccd1 vccd1 _16221_/D sky130_fd_sc_hd__clkbuf_1
X_10423_ _10428_/C vssd1 vssd1 vccd1 vccd1 _10440_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14191_ _14191_/A vssd1 vssd1 vccd1 vccd1 _16361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ _13423_/A vssd1 vssd1 vccd1 vccd1 _13364_/B sky130_fd_sc_hd__clkbuf_2
X_10354_ _15802_/Q _10362_/C _10204_/X vssd1 vssd1 vccd1 vccd1 _10354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _13073_/A vssd1 vssd1 vccd1 vccd1 _16202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10285_ _15789_/Q _10285_/B _10285_/C vssd1 vssd1 vccd1 vccd1 _10290_/A sky130_fd_sc_hd__and3_1
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12024_ _12059_/C vssd1 vssd1 vccd1 vccd1 _12065_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16674__79 vssd1 vssd1 vccd1 vccd1 _16674__79/HI _16750_/A sky130_fd_sc_hd__conb_1
XFILLER_93_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13975_ _13971_/Y _13973_/X _13974_/Y _13969_/C vssd1 vssd1 vccd1 vccd1 _13977_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_74_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15714_ _16551_/CLK _15714_/D vssd1 vssd1 vccd1 vccd1 _15714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _12963_/A _12926_/B _12926_/C vssd1 vssd1 vccd1 vccd1 _12927_/A sky130_fd_sc_hd__and3_1
X_16694_ _16694_/A _07792_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15645_ _15791_/CLK _15645_/D vssd1 vssd1 vccd1 vccd1 _15645_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _13705_/A vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__buf_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _16024_/Q _12031_/B _11814_/C vssd1 vssd1 vccd1 vccd1 _11810_/C sky130_fd_sc_hd__nand3_1
X_12788_ _12788_/A _12788_/B _12788_/C vssd1 vssd1 vccd1 vccd1 _12789_/A sky130_fd_sc_hd__and3_1
X_15576_ _16551_/CLK _15576_/D vssd1 vssd1 vccd1 vccd1 _15576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11739_ _11739_/A vssd1 vssd1 vccd1 vccd1 _16013_/D sky130_fd_sc_hd__clkbuf_1
X_14527_ _14535_/A _14527_/B _14527_/C vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__and3_1
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14458_ _16401_/Q _14458_/B _14458_/C vssd1 vssd1 vccd1 vccd1 _14458_/X sky130_fd_sc_hd__and3_1
XFILLER_128_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13409_ _16250_/Q _13467_/B _13416_/C vssd1 vssd1 vccd1 vccd1 _13409_/Y sky130_fd_sc_hd__nand3_1
X_14389_ _14555_/A _14389_/B _14389_/C vssd1 vssd1 vccd1 vccd1 _14390_/C sky130_fd_sc_hd__or3_1
XFILLER_143_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16128_ _16554_/Q _16128_/D vssd1 vssd1 vccd1 vccd1 _16128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08950_ _08950_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08951_/B sky130_fd_sc_hd__nor2_1
XFILLER_143_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16059_ _16118_/CLK _16059_/D vssd1 vssd1 vccd1 vccd1 _16059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07901_ _15660_/Q vssd1 vssd1 vccd1 vccd1 _09541_/C sky130_fd_sc_hd__clkinv_4
XFILLER_97_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08881_ _08706_/X _08879_/A _08833_/X vssd1 vssd1 vccd1 vccd1 _08882_/B sky130_fd_sc_hd__o21ai_1
XFILLER_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07832_ _07836_/A vssd1 vssd1 vccd1 vccd1 _07832_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07763_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__buf_12
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09502_ _09588_/A _09502_/B _09502_/C vssd1 vssd1 vccd1 vccd1 _09503_/A sky130_fd_sc_hd__and3_1
XFILLER_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09433_ _09427_/Y _09430_/X _09432_/Y vssd1 vssd1 vccd1 vccd1 _15620_/D sky130_fd_sc_hd__o21a_1
XFILLER_25_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _15611_/Q _09364_/B _09371_/C vssd1 vssd1 vccd1 vccd1 _09366_/C sky130_fd_sc_hd__nand3_1
XFILLER_80_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08315_ _08306_/A _08306_/B _08314_/Y vssd1 vssd1 vccd1 vccd1 _08414_/A sky130_fd_sc_hd__a21bo_1
X_09295_ _15355_/A _09295_/B vssd1 vssd1 vccd1 vccd1 _09296_/B sky130_fd_sc_hd__and2_1
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_20 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 _10729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_42 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08246_ _14785_/A _08066_/B _08245_/X vssd1 vssd1 vccd1 vccd1 _08253_/A sky130_fd_sc_hd__o21a_2
X_08177_ _08329_/B _08177_/B vssd1 vssd1 vccd1 vccd1 _08194_/A sky130_fd_sc_hd__and2_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10070_ _10697_/A vssd1 vssd1 vccd1 vccd1 _10578_/A sky130_fd_sc_hd__buf_2
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13760_ _16299_/Q _13760_/B _13765_/C vssd1 vssd1 vccd1 vccd1 _13760_/Y sky130_fd_sc_hd__nand3_1
X_10972_ _10970_/Y _10966_/C _10968_/Y _10969_/X vssd1 vssd1 vccd1 vccd1 _10973_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ _16152_/Q _12718_/C _12598_/X vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__a21o_1
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13691_ _14814_/A vssd1 vssd1 vccd1 vccd1 _13914_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12642_ _12924_/A vssd1 vssd1 vccd1 vccd1 _12868_/A sky130_fd_sc_hd__clkbuf_2
X_15430_ _16283_/Q _16285_/Q _16284_/Q _15428_/X vssd1 vssd1 vccd1 vccd1 _16606_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15361_ _09308_/X _15360_/A _09436_/A vssd1 vssd1 vccd1 vccd1 _15361_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12573_ _12653_/A _12573_/B _12580_/B vssd1 vssd1 vccd1 vccd1 _16131_/D sky130_fd_sc_hd__nor3_1
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11524_ _11525_/B _11525_/C _11525_/A vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__a21o_1
X_14312_ _14309_/Y _14310_/X _14311_/Y _14306_/C vssd1 vssd1 vccd1 vccd1 _14314_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15292_ _15292_/A _15292_/B vssd1 vssd1 vccd1 vccd1 _15292_/X sky130_fd_sc_hd__and2_1
XFILLER_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14243_ _14806_/A vssd1 vssd1 vccd1 vccd1 _14464_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_11455_ _16568_/Q vssd1 vssd1 vccd1 vccd1 _11473_/C sky130_fd_sc_hd__inv_2
XFILLER_109_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10406_ _10429_/A _10406_/B _10410_/B vssd1 vssd1 vccd1 vccd1 _15809_/D sky130_fd_sc_hd__nor3_1
X_14174_ _14175_/B _14175_/C _14175_/A vssd1 vssd1 vccd1 vccd1 _14176_/B sky130_fd_sc_hd__a21o_1
X_11386_ _11617_/A _11391_/C vssd1 vssd1 vccd1 vccd1 _11386_/X sky130_fd_sc_hd__or2_1
X_13125_ _16211_/Q _13135_/C _12901_/X vssd1 vssd1 vccd1 vccd1 _13125_/Y sky130_fd_sc_hd__a21oi_1
X_10337_ _10337_/A _10337_/B _10337_/C vssd1 vssd1 vccd1 vccd1 _10338_/C sky130_fd_sc_hd__nand3_1
XFILLER_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13072_/A _13056_/B _13056_/C vssd1 vssd1 vccd1 vccd1 _13057_/A sky130_fd_sc_hd__and3_1
X_10268_ _10268_/A _10268_/B vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__or2_1
XFILLER_87_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ _12292_/A vssd1 vssd1 vccd1 vccd1 _12007_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10199_ _10195_/Y _10197_/X _10198_/Y _10193_/C vssd1 vssd1 vccd1 vccd1 _10201_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16746_ _16746_/A _07762_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13958_ _16329_/Q _14179_/B _13958_/C vssd1 vssd1 vccd1 vccd1 _13958_/X sky130_fd_sc_hd__and3_1
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12909_ _16180_/Q _12916_/C _12850_/X vssd1 vssd1 vccd1 vccd1 _12909_/Y sky130_fd_sc_hd__a21oi_1
X_13889_ _13923_/C vssd1 vssd1 vccd1 vccd1 _13929_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15628_ _15791_/CLK _15628_/D vssd1 vssd1 vccd1 vccd1 _15628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15559_ _16551_/CLK _15559_/D vssd1 vssd1 vccd1 vccd1 _15559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08100_ _08100_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08114_/B sky130_fd_sc_hd__xor2_4
XFILLER_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09080_ _09294_/A vssd1 vssd1 vccd1 vccd1 _09240_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08031_ _15813_/Q vssd1 vssd1 vccd1 vccd1 _10332_/C sky130_fd_sc_hd__inv_2
XFILLER_135_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09982_ _14615_/A vssd1 vssd1 vccd1 vccd1 _09982_/X sky130_fd_sc_hd__buf_2
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08933_ _15521_/Q _08948_/C _08843_/X vssd1 vssd1 vccd1 vccd1 _08935_/B sky130_fd_sc_hd__a21oi_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08864_ _08946_/A _08864_/B _08868_/B vssd1 vssd1 vccd1 vccd1 _15501_/D sky130_fd_sc_hd__nor3_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07815_ _07818_/A vssd1 vssd1 vccd1 vccd1 _07815_/Y sky130_fd_sc_hd__inv_2
X_08795_ _14954_/A vssd1 vssd1 vccd1 vccd1 _09207_/A sky130_fd_sc_hd__buf_4
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09416_ _15621_/Q _09416_/B _09416_/C vssd1 vssd1 vccd1 vccd1 _09422_/A sky130_fd_sc_hd__and3_1
X_09347_ _09436_/A _09347_/B vssd1 vssd1 vccd1 vccd1 _09347_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ _09278_/A vssd1 vssd1 vccd1 vccd1 _09698_/A sky130_fd_sc_hd__buf_2
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08229_ _12473_/A _08229_/B vssd1 vssd1 vccd1 vccd1 _08229_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _15944_/Q _11465_/B _11246_/C vssd1 vssd1 vccd1 vccd1 _11242_/C sky130_fd_sc_hd__nand3_1
XFILLER_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11171_ _11171_/A vssd1 vssd1 vccd1 vccd1 _15933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10122_ _10152_/C vssd1 vssd1 vccd1 vccd1 _10158_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10053_ _10050_/Y _10059_/A _10052_/Y _10048_/C vssd1 vssd1 vccd1 vccd1 _10055_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14930_ _16475_/Q _14940_/C _14872_/X vssd1 vssd1 vccd1 vccd1 _14930_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16644__49 vssd1 vssd1 vccd1 vccd1 _16644__49/HI _16720_/A sky130_fd_sc_hd__conb_1
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14861_ _14859_/Y _14860_/X _14855_/C _14856_/C vssd1 vssd1 vccd1 vccd1 _14863_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_36_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16600_ _16607_/CLK _16600_/D vssd1 vssd1 vccd1 vccd1 _16600_/Q sky130_fd_sc_hd__dfxtp_1
X_13812_ _13812_/A vssd1 vssd1 vccd1 vccd1 _16306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14792_ _16454_/Q _14800_/C _14567_/X vssd1 vssd1 vccd1 vccd1 _14795_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16531_ _16595_/CLK _16531_/D vssd1 vssd1 vccd1 vccd1 _16531_/Q sky130_fd_sc_hd__dfxtp_1
X_10955_ _15904_/Q _10963_/C _10898_/X vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13743_ _16298_/Q _13745_/C _13570_/X vssd1 vssd1 vccd1 vccd1 _13743_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16462_ input11/X _16462_/D vssd1 vssd1 vccd1 vccd1 _16462_/Q sky130_fd_sc_hd__dfxtp_1
X_10886_ _14954_/A _10886_/B _10886_/C vssd1 vssd1 vccd1 vccd1 _10887_/C sky130_fd_sc_hd__or3_1
X_13674_ input2/X vssd1 vssd1 vccd1 vccd1 _14799_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15413_ _16181_/Q _16180_/Q _16179_/Q _15409_/X vssd1 vssd1 vccd1 vccd1 _16593_/D
+ sky130_fd_sc_hd__o31a_1
X_12625_ _12625_/A _12625_/B _12625_/C vssd1 vssd1 vccd1 vccd1 _12626_/A sky130_fd_sc_hd__and3_1
X_16393_ input11/X _16393_/D vssd1 vssd1 vccd1 vccd1 _16393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12556_ _12554_/Y _12548_/C _12550_/Y _12553_/X vssd1 vssd1 vccd1 vccd1 _12557_/C
+ sky130_fd_sc_hd__a211o_1
X_15344_ _15344_/A _15344_/B _15348_/B vssd1 vssd1 vccd1 vccd1 _16546_/D sky130_fd_sc_hd__nor3_1
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ _11509_/B _11509_/C _11282_/X vssd1 vssd1 vccd1 vccd1 _11510_/B sky130_fd_sc_hd__o21ai_1
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15275_ _15338_/A _15275_/B _15275_/C vssd1 vssd1 vccd1 vccd1 _15276_/A sky130_fd_sc_hd__and3_1
X_12487_ _16121_/Q _12487_/B _12487_/C vssd1 vssd1 vccd1 vccd1 _12487_/X sky130_fd_sc_hd__and3_1
X_11438_ _11435_/Y _11446_/A _11437_/Y _11431_/C vssd1 vssd1 vccd1 vccd1 _11440_/B
+ sky130_fd_sc_hd__o211a_1
X_14226_ _16367_/Q _14268_/C _14060_/X vssd1 vssd1 vccd1 vccd1 _14228_/B sky130_fd_sc_hd__a21oi_1
X_14157_ _14157_/A _14157_/B vssd1 vssd1 vccd1 vccd1 _14162_/C sky130_fd_sc_hd__nor2_1
X_11369_ _11366_/Y _11367_/X _11368_/Y _11364_/C vssd1 vssd1 vccd1 vccd1 _11371_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _13131_/A _13108_/B _13108_/C vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__and3_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14088_ _14084_/Y _14085_/X _14087_/Y _14082_/C vssd1 vssd1 vccd1 vccd1 _14090_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _16596_/Q vssd1 vssd1 vccd1 vccd1 _13053_/C sky130_fd_sc_hd__inv_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08580_ input10/X vssd1 vssd1 vccd1 vccd1 _12655_/A sky130_fd_sc_hd__buf_6
XFILLER_93_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16729_ _16729_/A _07834_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09201_ _09240_/A _09204_/C vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__and2_1
X_09132_ _15551_/Q _15550_/Q _15549_/Q _09090_/X vssd1 vssd1 vccd1 vccd1 _15561_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_148_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09063_ _10447_/A vssd1 vssd1 vccd1 vccd1 _09063_/X sky130_fd_sc_hd__buf_2
X_08014_ _08218_/B _08014_/B vssd1 vssd1 vccd1 vccd1 _08214_/B sky130_fd_sc_hd__nand2_2
XFILLER_118_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09965_ _09962_/A _09961_/Y _09962_/B vssd1 vssd1 vccd1 vccd1 _09965_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_134_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08916_ _08916_/A _08921_/C vssd1 vssd1 vccd1 vccd1 _08916_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09896_ _09749_/X _09891_/B _09895_/Y vssd1 vssd1 vccd1 vccd1 _15712_/D sky130_fd_sc_hd__o21a_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08847_ _15504_/Q _08849_/C _08805_/X vssd1 vssd1 vccd1 vccd1 _08851_/B sky130_fd_sc_hd__a21o_1
XFILLER_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08778_ _15488_/Q _08779_/C _08777_/X vssd1 vssd1 vccd1 vccd1 _08780_/A sky130_fd_sc_hd__a21oi_1
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ _10740_/A vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10671_ _10685_/C vssd1 vssd1 vccd1 vccd1 _10701_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12410_ _12410_/A _12418_/B vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__or2_1
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ _13390_/A vssd1 vssd1 vccd1 vccd1 _16247_/D sky130_fd_sc_hd__clkbuf_1
X_12341_ _12338_/Y _12339_/X _12340_/Y _12335_/C vssd1 vssd1 vccd1 vccd1 _12343_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_139_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15060_ _15271_/A _15064_/C vssd1 vssd1 vccd1 vccd1 _15060_/X sky130_fd_sc_hd__or2_1
X_12272_ _12268_/Y _12270_/X _12271_/Y _12266_/C vssd1 vssd1 vccd1 vccd1 _12274_/B
+ sky130_fd_sc_hd__o211ai_1
X_14011_ _14012_/B _14012_/C _14012_/A vssd1 vssd1 vccd1 vccd1 _14013_/B sky130_fd_sc_hd__a21o_1
X_11223_ _11334_/A vssd1 vssd1 vccd1 vccd1 _11264_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ _11151_/Y _11163_/A _11153_/Y _11148_/C vssd1 vssd1 vccd1 vccd1 _11156_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10105_ _15758_/Q _10106_/C _10104_/X vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__a21oi_1
X_15962_ _16005_/CLK _15962_/D vssd1 vssd1 vccd1 vccd1 _15962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11085_ _15922_/Q _11205_/B _11093_/C vssd1 vssd1 vccd1 vccd1 _11085_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10036_ _10036_/A vssd1 vssd1 vccd1 vccd1 _15743_/D sky130_fd_sc_hd__clkbuf_1
X_14913_ _14914_/B _14914_/C _14914_/A vssd1 vssd1 vccd1 vccd1 _14915_/B sky130_fd_sc_hd__a21o_1
X_15893_ _16553_/Q _15893_/D vssd1 vssd1 vccd1 vccd1 _15893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14844_ _14860_/C vssd1 vssd1 vccd1 vccd1 _14867_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14775_ _15005_/A _14780_/C vssd1 vssd1 vccd1 vccd1 _14775_/X sky130_fd_sc_hd__or2_1
X_11987_ _16049_/Q _12160_/B _11987_/C vssd1 vssd1 vccd1 vccd1 _11987_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16514_ _16607_/CLK _16514_/D vssd1 vssd1 vccd1 vccd1 _16514_/Q sky130_fd_sc_hd__dfxtp_1
X_13726_ _16295_/Q _13948_/B _13738_/C vssd1 vssd1 vccd1 vccd1 _13733_/A sky130_fd_sc_hd__and3_1
X_10938_ _11049_/A _10944_/C vssd1 vssd1 vccd1 vccd1 _10938_/X sky130_fd_sc_hd__or2_1
X_16445_ input11/X _16445_/D vssd1 vssd1 vccd1 vccd1 _16445_/Q sky130_fd_sc_hd__dfxtp_1
X_10869_ _15891_/Q _10929_/B _10878_/C vssd1 vssd1 vccd1 vccd1 _10869_/Y sky130_fd_sc_hd__nand3_1
X_13657_ _13696_/A _13657_/B _13657_/C vssd1 vssd1 vccd1 vccd1 _13658_/A sky130_fd_sc_hd__and3_1
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _12606_/Y _12607_/X _12602_/C _12603_/C vssd1 vssd1 vccd1 vccd1 _12610_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _16389_/CLK _16376_/D vssd1 vssd1 vccd1 vccd1 _16376_/Q sky130_fd_sc_hd__dfxtp_1
X_13588_ _13585_/Y _13594_/A _13587_/Y _13583_/C vssd1 vssd1 vccd1 vccd1 _13590_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15327_ _15327_/A _15327_/B vssd1 vssd1 vccd1 vccd1 _15327_/X sky130_fd_sc_hd__or2_1
X_12539_ _12540_/B _12540_/C _12540_/A vssd1 vssd1 vccd1 vccd1 _12541_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15258_ _15258_/A _15258_/B _15258_/C vssd1 vssd1 vccd1 vccd1 _15259_/A sky130_fd_sc_hd__and3_1
X_14209_ _14209_/A _14209_/B vssd1 vssd1 vccd1 vccd1 _14211_/B sky130_fd_sc_hd__nor2_1
X_15189_ _15187_/Y _15188_/X _15184_/C _15185_/C vssd1 vssd1 vccd1 vccd1 _15191_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_113_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ _09750_/A vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__clkbuf_2
X_08701_ _08630_/X _08690_/B _08694_/B _08700_/Y vssd1 vssd1 vccd1 vccd1 _15467_/D
+ sky130_fd_sc_hd__o31a_1
X_09681_ _09674_/C _09675_/C _09677_/Y _09687_/A vssd1 vssd1 vccd1 vccd1 _09687_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_55_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08632_ _10618_/A vssd1 vssd1 vccd1 vccd1 _08700_/A sky130_fd_sc_hd__buf_2
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08563_ _08555_/Y _08549_/Y _08562_/Y _08548_/B vssd1 vssd1 vccd1 vccd1 _08566_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _08494_/A _08446_/A vssd1 vssd1 vccd1 vccd1 _08494_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09115_ _09849_/A _09115_/B vssd1 vssd1 vccd1 vccd1 _09115_/X sky130_fd_sc_hd__or2_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09046_ _08883_/X _09044_/A _09045_/Y vssd1 vssd1 vccd1 vccd1 _15542_/D sky130_fd_sc_hd__o21a_1
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09948_ _15728_/Q _09992_/B _09955_/C vssd1 vssd1 vccd1 vccd1 _09950_/C sky130_fd_sc_hd__nand3_1
XFILLER_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09879_ _09879_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09879_/Y sky130_fd_sc_hd__nor2_1
X_11910_ _11930_/C vssd1 vssd1 vccd1 vccd1 _11944_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12890_ _12888_/Y _12889_/X _12883_/C _12884_/C vssd1 vssd1 vccd1 vccd1 _12892_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11948_/A _11841_/B _11845_/B vssd1 vssd1 vccd1 vccd1 _16027_/D sky130_fd_sc_hd__nor3_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _16019_/Q _11936_/B _11779_/C vssd1 vssd1 vccd1 vccd1 _11772_/X sky130_fd_sc_hd__and3_1
X_14560_ _14576_/C vssd1 vssd1 vccd1 vccd1 _14583_/C sky130_fd_sc_hd__clkbuf_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13511_/A vssd1 vssd1 vccd1 vccd1 _16264_/D sky130_fd_sc_hd__clkbuf_1
X_10723_ _10735_/C vssd1 vssd1 vccd1 vccd1 _10749_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _14720_/A _14496_/C vssd1 vssd1 vccd1 vccd1 _14491_/X sky130_fd_sc_hd__or2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _16261_/CLK _16230_/D vssd1 vssd1 vccd1 vccd1 _16230_/Q sky130_fd_sc_hd__dfxtp_2
X_13442_ _13498_/A _13442_/B _13447_/A vssd1 vssd1 vccd1 vccd1 _16254_/D sky130_fd_sc_hd__nor3_1
X_10654_ _10651_/Y _10660_/A _10653_/Y _10649_/C vssd1 vssd1 vccd1 vccd1 _10656_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16161_ _16237_/CLK _16161_/D vssd1 vssd1 vccd1 vccd1 _16161_/Q sky130_fd_sc_hd__dfxtp_1
X_13373_ _13374_/B _13374_/C _13264_/X vssd1 vssd1 vccd1 vccd1 _13375_/B sky130_fd_sc_hd__o21ai_1
X_10585_ _15844_/Q _10593_/C _10432_/X vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__a21o_1
XFILLER_139_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15112_ _15112_/A _15112_/B vssd1 vssd1 vccd1 vccd1 _15117_/C sky130_fd_sc_hd__nor2_1
XFILLER_126_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12324_ _16097_/Q _12332_/C _12323_/X vssd1 vssd1 vccd1 vccd1 _12324_/Y sky130_fd_sc_hd__a21oi_1
X_16092_ _16554_/Q _16092_/D vssd1 vssd1 vccd1 vccd1 _16092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15043_ _15040_/Y _15041_/X _15042_/Y _15038_/C vssd1 vssd1 vccd1 vccd1 _15045_/B
+ sky130_fd_sc_hd__o211ai_1
X_12255_ _16088_/Q _12318_/B _12263_/C vssd1 vssd1 vccd1 vccd1 _12257_/C sky130_fd_sc_hd__nand3_1
XFILLER_107_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11206_ _11203_/Y _11204_/X _11205_/Y _11200_/C vssd1 vssd1 vccd1 vccd1 _11208_/B
+ sky130_fd_sc_hd__o211ai_1
X_12186_ _12187_/B _12187_/C _12133_/X vssd1 vssd1 vccd1 vccd1 _12188_/B sky130_fd_sc_hd__o21ai_1
XFILLER_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11137_ _15929_/Q _11309_/B _11137_/C vssd1 vssd1 vccd1 vccd1 _11137_/Y sky130_fd_sc_hd__nand3_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15945_ _15365_/A _15945_/D vssd1 vssd1 vccd1 vccd1 _15945_/Q sky130_fd_sc_hd__dfxtp_1
X_11068_ _11068_/A vssd1 vssd1 vccd1 vccd1 _15919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10019_ _09307_/X _10017_/B _10012_/X vssd1 vssd1 vccd1 vccd1 _10019_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15876_ _16570_/CLK _15876_/D vssd1 vssd1 vccd1 vccd1 _15876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14827_ _14909_/A _14827_/B _14833_/B vssd1 vssd1 vccd1 vccd1 _16457_/D sky130_fd_sc_hd__nor3_1
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14758_ _14755_/Y _14756_/X _14757_/Y _14753_/C vssd1 vssd1 vccd1 vccd1 _14760_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_17_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13709_ _16293_/Q _13929_/B _13709_/C vssd1 vssd1 vccd1 vccd1 _13717_/B sky130_fd_sc_hd__and3_1
XFILLER_60_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14689_ _16437_/Q _14742_/B _14689_/C vssd1 vssd1 vccd1 vccd1 _14689_/X sky130_fd_sc_hd__and3_1
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16428_ _16607_/CLK _16428_/D vssd1 vssd1 vccd1 vccd1 _16428_/Q sky130_fd_sc_hd__dfxtp_1
X_16359_ _16389_/CLK _16359_/D vssd1 vssd1 vccd1 vccd1 _16359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09802_ _15699_/Q _10178_/B _09802_/C vssd1 vssd1 vccd1 vccd1 _09809_/A sky130_fd_sc_hd__and3_1
X_07994_ _16565_/Q vssd1 vssd1 vccd1 vccd1 _11287_/A sky130_fd_sc_hd__inv_2
X_09733_ _09733_/A _09733_/B vssd1 vssd1 vccd1 vccd1 _09733_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09664_ _15659_/Q _15658_/Q _15657_/Q _09536_/X vssd1 vssd1 vccd1 vccd1 _15669_/D
+ sky130_fd_sc_hd__o31a_1
X_08615_ _10501_/A vssd1 vssd1 vccd1 vccd1 _15346_/B sky130_fd_sc_hd__buf_2
XFILLER_55_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09595_ _09595_/A _09595_/B _09598_/B vssd1 vssd1 vccd1 vccd1 _15654_/D sky130_fd_sc_hd__nor3_1
XFILLER_43_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _15452_/Q _08561_/B _15315_/C vssd1 vssd1 vccd1 vccd1 _08555_/A sky130_fd_sc_hd__a21o_1
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08477_ _08491_/B _08477_/B vssd1 vssd1 vccd1 vccd1 _08479_/B sky130_fd_sc_hd__xor2_1
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10370_ _10573_/A _10370_/B vssd1 vssd1 vccd1 vccd1 _10370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09029_ _09029_/A _09029_/B vssd1 vssd1 vccd1 vccd1 _09031_/A sky130_fd_sc_hd__or2_1
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12040_ _12033_/C _12034_/C _12037_/Y _12038_/X vssd1 vssd1 vccd1 vccd1 _12041_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13991_ _13991_/A _13991_/B vssd1 vssd1 vccd1 vccd1 _13992_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15730_ _15812_/CLK _15730_/D vssd1 vssd1 vccd1 vccd1 _15730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12942_ _12963_/A _12942_/B _12942_/C vssd1 vssd1 vccd1 vccd1 _12943_/A sky130_fd_sc_hd__and3_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15661_ _15791_/CLK _15661_/D vssd1 vssd1 vccd1 vccd1 _15661_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12873_ _12896_/C vssd1 vssd1 vccd1 vccd1 _12910_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14839_/A _14612_/B _14612_/C vssd1 vssd1 vccd1 vccd1 _14613_/C sky130_fd_sc_hd__or3_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _11832_/A _11824_/B _11824_/C vssd1 vssd1 vccd1 vccd1 _11825_/A sky130_fd_sc_hd__and3_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _16551_/CLK _15592_/D vssd1 vssd1 vccd1 vccd1 _15592_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _14624_/A _14543_/B _14549_/B vssd1 vssd1 vccd1 vccd1 _16412_/D sky130_fd_sc_hd__nor3_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _12605_/A vssd1 vssd1 vccd1 vccd1 _11755_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _15866_/Q _10707_/C _08748_/A vssd1 vssd1 vccd1 vccd1 _10708_/A sky130_fd_sc_hd__a21oi_1
X_14474_ _14471_/Y _14472_/X _14473_/Y _14469_/C vssd1 vssd1 vccd1 vccd1 _14476_/B
+ sky130_fd_sc_hd__o211ai_1
X_11686_ _11721_/C vssd1 vssd1 vccd1 vccd1 _11729_/C sky130_fd_sc_hd__clkbuf_2
X_16213_ _16237_/CLK _16213_/D vssd1 vssd1 vccd1 vccd1 _16213_/Q sky130_fd_sc_hd__dfxtp_1
X_13425_ _13425_/A _13432_/B vssd1 vssd1 vccd1 vccd1 _13427_/A sky130_fd_sc_hd__or2_1
X_10637_ _10637_/A vssd1 vssd1 vccd1 vccd1 _15851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16144_ _16261_/CLK _16144_/D vssd1 vssd1 vccd1 vccd1 _16144_/Q sky130_fd_sc_hd__dfxtp_1
X_10568_ _11384_/A vssd1 vssd1 vccd1 vccd1 _10759_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13356_ _16244_/Q _13364_/C _13133_/X vssd1 vssd1 vccd1 vccd1 _13356_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12307_ _12307_/A vssd1 vssd1 vccd1 vccd1 _12325_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16075_ _16118_/CLK _16075_/D vssd1 vssd1 vccd1 vccd1 _16075_/Q sky130_fd_sc_hd__dfxtp_1
X_13287_ _13287_/A vssd1 vssd1 vccd1 vccd1 _16232_/D sky130_fd_sc_hd__clkbuf_1
X_10499_ _10740_/A vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15026_ _16491_/Q _15035_/C _14858_/X vssd1 vssd1 vccd1 vccd1 _15026_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12238_ _12236_/A _12236_/B _12237_/X vssd1 vssd1 vccd1 vccd1 _16084_/D sky130_fd_sc_hd__a21oi_1
XFILLER_111_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12169_ _12167_/Y _12163_/C _12165_/Y _12166_/X vssd1 vssd1 vccd1 vccd1 _12170_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_6
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15928_ _16005_/CLK _15928_/D vssd1 vssd1 vccd1 vccd1 _15928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15859_ _16595_/CLK _15859_/D vssd1 vssd1 vccd1 vccd1 _15859_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08400_ _08400_/A _08400_/B vssd1 vssd1 vccd1 vccd1 _08400_/Y sky130_fd_sc_hd__nor2_1
X_09380_ _09378_/A _09378_/B _09377_/Y _09379_/Y vssd1 vssd1 vccd1 vccd1 _15610_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08331_ _08331_/A _08160_/A vssd1 vssd1 vccd1 vccd1 _08336_/B sky130_fd_sc_hd__or2b_1
XFILLER_33_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08262_ _15462_/Q vssd1 vssd1 vccd1 vccd1 _15335_/C sky130_fd_sc_hd__clkinv_2
X_08193_ _08346_/A _08346_/B vssd1 vssd1 vccd1 vccd1 _08194_/B sky130_fd_sc_hd__xor2_4
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07977_ _16611_/Q vssd1 vssd1 vccd1 vccd1 _13886_/A sky130_fd_sc_hd__clkinv_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09716_ _09801_/A vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09647_ _09643_/A _09642_/Y _09643_/B vssd1 vssd1 vccd1 vccd1 _09647_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_35_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09581_/C vssd1 vssd1 vccd1 vccd1 _09592_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08529_/A _08529_/B vssd1 vssd1 vccd1 vccd1 _08530_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ _11540_/A vssd1 vssd1 vccd1 vccd1 _15985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11471_ _12605_/A vssd1 vssd1 vccd1 vccd1 _11471_/X sky130_fd_sc_hd__clkbuf_2
X_10422_ _15831_/Q vssd1 vssd1 vccd1 vccd1 _10428_/C sky130_fd_sc_hd__inv_2
X_13210_ _13246_/A _13210_/B _13210_/C vssd1 vssd1 vccd1 vccd1 _13211_/A sky130_fd_sc_hd__and3_1
X_14190_ _14197_/A _14190_/B _14190_/C vssd1 vssd1 vccd1 vccd1 _14191_/A sky130_fd_sc_hd__and3_1
X_10353_ _10353_/A vssd1 vssd1 vccd1 vccd1 _15799_/D sky130_fd_sc_hd__clkbuf_1
X_13141_ _16213_/Q _13143_/C _13140_/X vssd1 vssd1 vccd1 vccd1 _13144_/A sky130_fd_sc_hd__a21oi_1
XFILLER_124_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13072_ _13072_/A _13072_/B _13072_/C vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__and3_1
XFILLER_3_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10284_ _15789_/Q _10313_/B _10176_/X vssd1 vssd1 vccd1 vccd1 _10286_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12023_ _12045_/C vssd1 vssd1 vccd1 vccd1 _12059_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13974_ _16330_/Q _14032_/B _13981_/C vssd1 vssd1 vccd1 vccd1 _13974_/Y sky130_fd_sc_hd__nand3_1
X_15713_ _15812_/CLK _15713_/D vssd1 vssd1 vccd1 vccd1 _15713_/Q sky130_fd_sc_hd__dfxtp_1
X_12925_ _13151_/A _12925_/B _12925_/C vssd1 vssd1 vccd1 vccd1 _12926_/C sky130_fd_sc_hd__or3_1
X_16693_ _16693_/A _07791_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15644_ _15791_/CLK _15644_/D vssd1 vssd1 vccd1 vccd1 _15644_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12856_ _12936_/A _12856_/B _12862_/B vssd1 vssd1 vccd1 vccd1 _16171_/D sky130_fd_sc_hd__nor3_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _12373_/A vssd1 vssd1 vccd1 vccd1 _12031_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _16551_/CLK _15575_/D vssd1 vssd1 vccd1 vccd1 _15575_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12785_/Y _12781_/C _12783_/Y _12784_/X vssd1 vssd1 vccd1 vccd1 _12788_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_42_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14524_/Y _14519_/C _14521_/Y _14523_/X vssd1 vssd1 vccd1 vccd1 _14527_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_14_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11738_ _11776_/A _11738_/B _11738_/C vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__and3_1
XFILLER_30_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14457_ _16401_/Q _14466_/C _14294_/X vssd1 vssd1 vccd1 vccd1 _14457_/Y sky130_fd_sc_hd__a21oi_1
X_11669_ _11669_/A _11679_/B vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__or2_1
XFILLER_128_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13408_ _16251_/Q _13631_/B _13416_/C vssd1 vssd1 vccd1 vccd1 _13408_/X sky130_fd_sc_hd__and3_1
X_14388_ _14389_/B _14389_/C _14387_/X vssd1 vssd1 vccd1 vccd1 _14390_/B sky130_fd_sc_hd__o21ai_1
XFILLER_128_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16127_ _16554_/Q _16127_/D vssd1 vssd1 vccd1 vccd1 _16127_/Q sky130_fd_sc_hd__dfxtp_1
X_13339_ _13354_/A _13339_/B _13339_/C vssd1 vssd1 vccd1 vccd1 _13340_/A sky130_fd_sc_hd__and3_1
XFILLER_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16058_ _16118_/CLK _16058_/D vssd1 vssd1 vccd1 vccd1 _16058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07900_ _08295_/A _07900_/B vssd1 vssd1 vccd1 vccd1 _08100_/A sky130_fd_sc_hd__xnor2_4
X_15009_ _15117_/A _15009_/B _15009_/C vssd1 vssd1 vccd1 vccd1 _15010_/C sky130_fd_sc_hd__or3_1
X_08880_ _08921_/A _08921_/B _08880_/C vssd1 vssd1 vccd1 vccd1 _08882_/A sky130_fd_sc_hd__and3_1
X_07831_ _07837_/A vssd1 vssd1 vccd1 vccd1 _07836_/A sky130_fd_sc_hd__buf_12
XFILLER_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07762_ _07762_/A vssd1 vssd1 vccd1 vccd1 _07762_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09501_ _09501_/A _09501_/B _09501_/C vssd1 vssd1 vccd1 vccd1 _09502_/C sky130_fd_sc_hd__nand3_1
XFILLER_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09432_ _09427_/Y _09430_/X _09431_/X vssd1 vssd1 vccd1 vccd1 _09432_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09363_ _15611_/Q _09371_/C _09362_/X vssd1 vssd1 vccd1 vccd1 _09366_/B sky130_fd_sc_hd__a21o_1
X_08314_ _08314_/A _08314_/B vssd1 vssd1 vccd1 vccd1 _08314_/Y sky130_fd_sc_hd__nand2_1
X_09294_ _09294_/A vssd1 vssd1 vccd1 vccd1 _15355_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_10 _10060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_32 _11150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 _10285_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ _08245_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08245_/X sky130_fd_sc_hd__or2_1
XFILLER_21_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08176_ _08176_/A _08176_/B vssd1 vssd1 vccd1 vccd1 _08177_/B sky130_fd_sc_hd__or2_1
XFILLER_119_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10971_ _10968_/Y _10969_/X _10970_/Y _10966_/C vssd1 vssd1 vccd1 vccd1 _10973_/B
+ sky130_fd_sc_hd__o211ai_1
X_12710_ _12796_/A _12710_/B _12714_/A vssd1 vssd1 vccd1 vccd1 _16150_/D sky130_fd_sc_hd__nor3_1
XFILLER_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13690_ input4/X vssd1 vssd1 vccd1 vccd1 _14814_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12641_ _12643_/B _12643_/C _12416_/X vssd1 vssd1 vccd1 vccd1 _12644_/B sky130_fd_sc_hd__o21ai_1
X_15360_ _15360_/A _15360_/B vssd1 vssd1 vccd1 vccd1 _16550_/D sky130_fd_sc_hd__nor2_1
X_12572_ _12570_/Y _12565_/C _12568_/Y _12580_/A vssd1 vssd1 vccd1 vccd1 _12580_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_8_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14311_ _16378_/Q _14311_/B _14317_/C vssd1 vssd1 vccd1 vccd1 _14311_/Y sky130_fd_sc_hd__nand3_1
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11523_ _15984_/Q _11750_/B _11529_/C vssd1 vssd1 vccd1 vccd1 _11525_/C sky130_fd_sc_hd__nand3_1
X_15291_ _15291_/A _15291_/B vssd1 vssd1 vccd1 vccd1 _15292_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14242_ _16370_/Q _14245_/C _14132_/X vssd1 vssd1 vccd1 vccd1 _14242_/Y sky130_fd_sc_hd__a21oi_1
X_11454_ _11454_/A vssd1 vssd1 vccd1 vccd1 _15973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ _10403_/Y _10399_/C _10401_/Y _10410_/A vssd1 vssd1 vccd1 vccd1 _10410_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11385_ _11385_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11391_/C sky130_fd_sc_hd__nor2_1
X_14173_ _16360_/Q _14289_/B _14179_/C vssd1 vssd1 vccd1 vccd1 _14175_/C sky130_fd_sc_hd__nand3_1
XFILLER_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124_ _13124_/A vssd1 vssd1 vccd1 vccd1 _16209_/D sky130_fd_sc_hd__clkbuf_1
X_10336_ _10337_/B _10337_/C _10337_/A vssd1 vssd1 vccd1 vccd1 _10338_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _15785_/Q _10463_/B _10267_/C vssd1 vssd1 vccd1 vccd1 _10268_/B sky130_fd_sc_hd__and3_1
X_13055_ _13049_/C _13050_/C _13052_/Y _13053_/X vssd1 vssd1 vccd1 vccd1 _13056_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12006_ _12084_/A _12006_/B _12012_/B vssd1 vssd1 vccd1 vccd1 _16051_/D sky130_fd_sc_hd__nor3_1
X_10198_ _15773_/Q _10396_/B _10206_/C vssd1 vssd1 vccd1 vccd1 _10198_/Y sky130_fd_sc_hd__nand3_1
XFILLER_120_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16745_ _16745_/A _07761_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
XFILLER_81_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13957_ _14799_/A vssd1 vssd1 vccd1 vccd1 _14179_/B sky130_fd_sc_hd__clkbuf_2
X_12908_ _12908_/A vssd1 vssd1 vccd1 vccd1 _16178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13888_ _13908_/C vssd1 vssd1 vccd1 vccd1 _13923_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15627_ _15791_/CLK _15627_/D vssd1 vssd1 vccd1 vccd1 _15627_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ _12847_/A _12839_/B _12839_/C vssd1 vssd1 vccd1 vccd1 _12840_/A sky130_fd_sc_hd__and3_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15558_ _16551_/CLK _15558_/D vssd1 vssd1 vccd1 vccd1 _15558_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14509_ _16409_/Q _14569_/B _14516_/C vssd1 vssd1 vccd1 vccd1 _14511_/C sky130_fd_sc_hd__nand3_1
X_15489_ _16570_/CLK _15489_/D vssd1 vssd1 vccd1 vccd1 _15489_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08030_ _16415_/Q vssd1 vssd1 vccd1 vccd1 _14444_/A sky130_fd_sc_hd__inv_2
XFILLER_128_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09981_ _15415_/A vssd1 vssd1 vccd1 vccd1 _14615_/A sky130_fd_sc_hd__buf_2
XFILLER_131_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08932_ _08937_/C vssd1 vssd1 vccd1 vccd1 _08948_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_97_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08863_ _08851_/C _08852_/C _08860_/Y _08868_/A vssd1 vssd1 vccd1 vccd1 _08868_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07814_ _07818_/A vssd1 vssd1 vccd1 vccd1 _07814_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08794_ _14895_/A vssd1 vssd1 vccd1 vccd1 _14954_/A sky130_fd_sc_hd__buf_2
XFILLER_38_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09415_ _15621_/Q _09416_/C _09369_/X vssd1 vssd1 vccd1 vccd1 _09415_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09346_ _15355_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09347_/B sky130_fd_sc_hd__and2_1
XFILLER_139_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09277_ _09277_/A _09277_/B vssd1 vssd1 vccd1 vccd1 _09277_/X sky130_fd_sc_hd__or2_1
XFILLER_148_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08228_ _08228_/A vssd1 vssd1 vccd1 vccd1 _08228_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08159_ _08330_/A _08330_/B vssd1 vssd1 vccd1 vccd1 _08331_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ _11208_/A _11170_/B _11170_/C vssd1 vssd1 vccd1 vccd1 _11171_/A sky130_fd_sc_hd__and3_1
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10121_ _10133_/C vssd1 vssd1 vccd1 vccd1 _10152_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10052_ _15747_/Q _10308_/C _10057_/C vssd1 vssd1 vccd1 vccd1 _10052_/Y sky130_fd_sc_hd__nand3_1
XFILLER_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14860_ _16464_/Q _15027_/B _14860_/C vssd1 vssd1 vccd1 vccd1 _14860_/X sky130_fd_sc_hd__and3_1
XFILLER_75_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13811_ _13811_/A _13811_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _13812_/A sky130_fd_sc_hd__and3_1
X_14791_ _14909_/A _14791_/B _14795_/A vssd1 vssd1 vccd1 vccd1 _16452_/D sky130_fd_sc_hd__nor3_1
XFILLER_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16530_ _16595_/CLK _16530_/D vssd1 vssd1 vccd1 vccd1 _16530_/Q sky130_fd_sc_hd__dfxtp_1
X_13742_ _13742_/A vssd1 vssd1 vccd1 vccd1 _16296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10954_ _10954_/A _10954_/B _10959_/A vssd1 vssd1 vccd1 vccd1 _15902_/D sky130_fd_sc_hd__nor3_1
XFILLER_44_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16461_ input11/X _16461_/D vssd1 vssd1 vccd1 vccd1 _16461_/Q sky130_fd_sc_hd__dfxtp_2
X_13673_ _16289_/Q _13684_/C _13450_/X vssd1 vssd1 vccd1 vccd1 _13673_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10885_ _10886_/B _10886_/C _09978_/X vssd1 vssd1 vccd1 vccd1 _10887_/B sky130_fd_sc_hd__o21ai_1
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15412_ _16173_/Q _16172_/Q _16171_/Q _15409_/X vssd1 vssd1 vccd1 vccd1 _16592_/D
+ sky130_fd_sc_hd__o31a_1
X_12624_ _12622_/Y _12617_/C _12620_/Y _12621_/X vssd1 vssd1 vccd1 vccd1 _12625_/C
+ sky130_fd_sc_hd__a211o_1
X_16392_ input11/X _16392_/D vssd1 vssd1 vccd1 vccd1 _16392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15343_ _15337_/C _15338_/C _15340_/Y _15348_/A vssd1 vssd1 vccd1 vccd1 _15348_/B
+ sky130_fd_sc_hd__a211oi_1
X_12555_ _12550_/Y _12553_/X _12554_/Y _12548_/C vssd1 vssd1 vccd1 vccd1 _12557_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_12_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11506_ _11619_/A vssd1 vssd1 vccd1 vccd1 _11547_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15274_ _15274_/A _15274_/B _15274_/C vssd1 vssd1 vccd1 vccd1 _15275_/C sky130_fd_sc_hd__or3_1
X_12486_ _16121_/Q _12495_/C _12323_/X vssd1 vssd1 vccd1 vccd1 _12486_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14225_ _14260_/C vssd1 vssd1 vccd1 vccd1 _14268_/C sky130_fd_sc_hd__clkbuf_2
X_11437_ _15971_/Q _11495_/B _11444_/C vssd1 vssd1 vccd1 vccd1 _11437_/Y sky130_fd_sc_hd__nand3_1
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14156_ _14156_/A _14156_/B vssd1 vssd1 vccd1 vccd1 _14157_/B sky130_fd_sc_hd__nor2_1
X_11368_ _15962_/Q _11488_/B _11375_/C vssd1 vssd1 vccd1 vccd1 _11368_/Y sky130_fd_sc_hd__nand3_1
XFILLER_4_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13107_ _13107_/A _13107_/B _13107_/C vssd1 vssd1 vccd1 vccd1 _13108_/C sky130_fd_sc_hd__nand3_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _10521_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10319_/X sky130_fd_sc_hd__or2_1
XFILLER_140_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _16346_/Q _14311_/B _14094_/C vssd1 vssd1 vccd1 vccd1 _14087_/Y sky130_fd_sc_hd__nand3_1
X_11299_ _11299_/A vssd1 vssd1 vccd1 vccd1 _15951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13038_/A vssd1 vssd1 vccd1 vccd1 _16197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14989_ _16483_/Q _15149_/B _14995_/C vssd1 vssd1 vccd1 vccd1 _14989_/Y sky130_fd_sc_hd__nand3_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16728_ _16728_/A _07833_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09200_ _09076_/X _09193_/B _09196_/B _09199_/Y vssd1 vssd1 vccd1 vccd1 _15575_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_62_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09131_ _09087_/X _09128_/A _09130_/Y vssd1 vssd1 vccd1 vccd1 _15560_/D sky130_fd_sc_hd__o21a_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09062_ _09400_/A vssd1 vssd1 vccd1 vccd1 _09148_/A sky130_fd_sc_hd__clkbuf_2
X_08013_ _08218_/A _08012_/C _16559_/Q vssd1 vssd1 vccd1 vccd1 _08014_/B sky130_fd_sc_hd__a21o_1
XFILLER_116_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09964_ _09962_/A _09962_/B _09961_/Y _09963_/Y vssd1 vssd1 vccd1 vccd1 _15727_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08915_ _08908_/B _08912_/B _08914_/X vssd1 vssd1 vccd1 vccd1 _08921_/C sky130_fd_sc_hd__o21a_1
X_09895_ _09658_/X _09891_/B _09894_/X vssd1 vssd1 vccd1 vccd1 _09895_/Y sky130_fd_sc_hd__a21oi_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08846_ _08846_/A _08846_/B _08851_/A vssd1 vssd1 vccd1 vccd1 _15499_/D sky130_fd_sc_hd__nor3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ _15346_/B vssd1 vssd1 vccd1 vccd1 _08777_/X sky130_fd_sc_hd__buf_2
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10670_ _10675_/C vssd1 vssd1 vccd1 vccd1 _10685_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _15603_/Q _09416_/B _09329_/C vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__and3_1
X_12340_ _16098_/Q _12340_/B _12346_/C vssd1 vssd1 vccd1 vccd1 _12340_/Y sky130_fd_sc_hd__nand3_1
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12271_ _16089_/Q _12443_/B _12271_/C vssd1 vssd1 vccd1 vccd1 _12271_/Y sky130_fd_sc_hd__nand3_1
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _16336_/Q _14010_/B _14017_/C vssd1 vssd1 vccd1 vccd1 _14012_/C sky130_fd_sc_hd__nand3_1
X_11222_ _11220_/A _11220_/B _11221_/X vssd1 vssd1 vccd1 vccd1 _15940_/D sky130_fd_sc_hd__a21oi_1
XFILLER_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _15931_/Q _11212_/B _11161_/C vssd1 vssd1 vccd1 vccd1 _11153_/Y sky130_fd_sc_hd__nand3_1
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10104_ _10755_/B vssd1 vssd1 vccd1 vccd1 _10104_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15961_ _16005_/CLK _15961_/D vssd1 vssd1 vccd1 vccd1 _15961_/Q sky130_fd_sc_hd__dfxtp_1
X_11084_ _15923_/Q _11084_/B _11093_/C vssd1 vssd1 vccd1 vccd1 _11084_/X sky130_fd_sc_hd__and3_1
XFILLER_49_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10035_ _10082_/A _10035_/B _10035_/C vssd1 vssd1 vccd1 vccd1 _10036_/A sky130_fd_sc_hd__and3_1
X_14912_ _16472_/Q _15129_/B _14918_/C vssd1 vssd1 vccd1 vccd1 _14914_/C sky130_fd_sc_hd__nand3_1
XFILLER_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15892_ _16553_/Q _15892_/D vssd1 vssd1 vccd1 vccd1 _15892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14843_ _16478_/Q vssd1 vssd1 vccd1 vccd1 _14860_/C sky130_fd_sc_hd__inv_2
XFILLER_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ _14774_/A _14774_/B vssd1 vssd1 vccd1 vccd1 _14780_/C sky130_fd_sc_hd__nor2_1
X_11986_ _16050_/Q _12210_/B _11987_/C vssd1 vssd1 vccd1 vccd1 _11986_/X sky130_fd_sc_hd__and3_1
XFILLER_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16513_ _16607_/CLK _16513_/D vssd1 vssd1 vccd1 vccd1 _16513_/Q sky130_fd_sc_hd__dfxtp_1
X_13725_ _13725_/A vssd1 vssd1 vccd1 vccd1 _13948_/B sky130_fd_sc_hd__clkbuf_2
X_10937_ _10937_/A _10937_/B vssd1 vssd1 vccd1 vccd1 _10944_/C sky130_fd_sc_hd__nor2_1
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ _16607_/CLK _16444_/D vssd1 vssd1 vccd1 vccd1 _16444_/Q sky130_fd_sc_hd__dfxtp_1
X_13656_ _13717_/A _13656_/B _13656_/C vssd1 vssd1 vccd1 vccd1 _13657_/C sky130_fd_sc_hd__or3_1
X_10868_ _15892_/Q _11039_/B _10868_/C vssd1 vssd1 vccd1 vccd1 _10880_/A sky130_fd_sc_hd__and3_1
X_12607_ _16137_/Q _12770_/B _12607_/C vssd1 vssd1 vccd1 vccd1 _12607_/X sky130_fd_sc_hd__and3_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _16389_/CLK _16375_/D vssd1 vssd1 vccd1 vccd1 _16375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13587_ _16275_/Q _13760_/B _13592_/C vssd1 vssd1 vccd1 vccd1 _13587_/Y sky130_fd_sc_hd__nand3_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _10796_/Y _10797_/X _10798_/Y _10794_/C vssd1 vssd1 vccd1 vccd1 _10801_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_40_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15326_ _15366_/B _15326_/B _15325_/X vssd1 vssd1 vccd1 vccd1 _16541_/D sky130_fd_sc_hd__nor3b_1
XFILLER_118_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12538_ _16128_/Q _12600_/B _12545_/C vssd1 vssd1 vccd1 vccd1 _12540_/C sky130_fd_sc_hd__nand3_1
X_15257_ _15255_/Y _15251_/C _15253_/Y _15254_/X vssd1 vssd1 vccd1 vccd1 _15258_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12469_ _12470_/B _12470_/C _12416_/X vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__o21ai_1
XFILLER_99_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14208_ _14208_/A _14217_/B vssd1 vssd1 vccd1 vccd1 _14211_/A sky130_fd_sc_hd__or2_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15188_ _16518_/Q _15241_/B _15188_/C vssd1 vssd1 vccd1 vccd1 _15188_/X sky130_fd_sc_hd__and3_1
XFILLER_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14139_ _14139_/A vssd1 vssd1 vccd1 vccd1 _16353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08700_ _08700_/A _08705_/C vssd1 vssd1 vccd1 vccd1 _08700_/Y sky130_fd_sc_hd__nor2_1
X_09680_ _09677_/Y _09687_/A _09674_/C _09675_/C vssd1 vssd1 vccd1 vccd1 _09682_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08631_ _09278_/A vssd1 vssd1 vccd1 vccd1 _10618_/A sky130_fd_sc_hd__buf_2
XFILLER_82_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08562_ _15327_/A _08568_/B vssd1 vssd1 vccd1 vccd1 _08562_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08493_ _08475_/A _08475_/B _08492_/X vssd1 vssd1 vccd1 vccd1 _08534_/B sky130_fd_sc_hd__o21ai_2
XFILLER_120_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09114_ _09114_/A _09114_/B vssd1 vssd1 vccd1 vccd1 _09115_/B sky130_fd_sc_hd__nor2_1
X_09045_ _09006_/X _09044_/A _08927_/X vssd1 vssd1 vccd1 vccd1 _09045_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09947_ _15728_/Q _09955_/C _08589_/A vssd1 vssd1 vccd1 vccd1 _09950_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09878_ _15712_/Q _09919_/B _09884_/C vssd1 vssd1 vccd1 vccd1 _09880_/B sky130_fd_sc_hd__and3_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08829_ _08916_/A _08836_/C vssd1 vssd1 vccd1 vccd1 _08829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11838_/Y _11832_/C _11835_/Y _11845_/A vssd1 vssd1 vccd1 vccd1 _11845_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _16019_/Q _11779_/C _11770_/X vssd1 vssd1 vccd1 vccd1 _11771_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13510_ _13526_/A _13510_/B _13510_/C vssd1 vssd1 vccd1 vccd1 _13511_/A sky130_fd_sc_hd__and3_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10722_ _10726_/C vssd1 vssd1 vccd1 vccd1 _10735_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _14490_/A _14490_/B vssd1 vssd1 vccd1 vccd1 _14496_/C sky130_fd_sc_hd__nor2_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ _16255_/Q _13665_/B _13452_/C vssd1 vssd1 vccd1 vccd1 _13447_/A sky130_fd_sc_hd__and3_1
XFILLER_41_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10653_ _15855_/Q _10702_/B _10658_/C vssd1 vssd1 vccd1 vccd1 _10653_/Y sky130_fd_sc_hd__nand3_1
XFILLER_139_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16160_ _16261_/CLK _16160_/D vssd1 vssd1 vccd1 vccd1 _16160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13372_ _13598_/A vssd1 vssd1 vccd1 vccd1 _13412_/A sky130_fd_sc_hd__clkbuf_2
X_10584_ _10676_/A _10584_/B _10588_/A vssd1 vssd1 vccd1 vccd1 _15841_/D sky130_fd_sc_hd__nor3_1
X_15111_ _15111_/A _15111_/B vssd1 vssd1 vccd1 vccd1 _15112_/B sky130_fd_sc_hd__nor2_1
X_12323_ _12605_/A vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__clkbuf_2
X_16091_ _16118_/CLK _16091_/D vssd1 vssd1 vccd1 vccd1 _16091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15042_ _16492_/Q _15149_/B _15049_/C vssd1 vssd1 vccd1 vccd1 _15042_/Y sky130_fd_sc_hd__nand3_1
XFILLER_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12254_ _16088_/Q _12263_/C _12029_/X vssd1 vssd1 vccd1 vccd1 _12257_/B sky130_fd_sc_hd__a21o_1
XFILLER_141_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11205_ _15938_/Q _11205_/B _11211_/C vssd1 vssd1 vccd1 vccd1 _11205_/Y sky130_fd_sc_hd__nand3_1
XFILLER_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12185_ _12185_/A vssd1 vssd1 vccd1 vccd1 _12222_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11136_ _15930_/Q _11359_/B _11137_/C vssd1 vssd1 vccd1 vccd1 _11136_/X sky130_fd_sc_hd__and3_1
XFILLER_110_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15944_ _15365_/A _15944_/D vssd1 vssd1 vccd1 vccd1 _15944_/Q sky130_fd_sc_hd__dfxtp_1
X_11067_ _11088_/A _11067_/B _11067_/C vssd1 vssd1 vccd1 vccd1 _11068_/A sky130_fd_sc_hd__and3_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10018_ _08644_/X _10016_/B _10017_/Y vssd1 vssd1 vccd1 vccd1 _15738_/D sky130_fd_sc_hd__o21a_1
X_15875_ _16570_/CLK _15875_/D vssd1 vssd1 vccd1 vccd1 _15875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14826_ _14824_/Y _14819_/C _14822_/Y _14833_/A vssd1 vssd1 vccd1 vccd1 _14833_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_45_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14757_ _16447_/Q _14875_/B _14764_/C vssd1 vssd1 vccd1 vccd1 _14757_/Y sky130_fd_sc_hd__nand3_1
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11969_ _16047_/Q _11969_/B _11979_/C vssd1 vssd1 vccd1 vccd1 _11974_/A sky130_fd_sc_hd__and3_1
XFILLER_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13708_ _14830_/A vssd1 vssd1 vccd1 vccd1 _13929_/B sky130_fd_sc_hd__clkbuf_2
X_14688_ _16437_/Q _14697_/C _14574_/X vssd1 vssd1 vccd1 vccd1 _14688_/Y sky130_fd_sc_hd__a21oi_1
X_16427_ _16607_/CLK _16427_/D vssd1 vssd1 vccd1 vccd1 _16427_/Q sky130_fd_sc_hd__dfxtp_1
X_13639_ _16284_/Q _13869_/B _13639_/C vssd1 vssd1 vccd1 vccd1 _13647_/A sky130_fd_sc_hd__and3_1
X_16358_ _16389_/CLK _16358_/D vssd1 vssd1 vccd1 vccd1 _16358_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15309_ _15324_/A _15309_/B vssd1 vssd1 vccd1 vccd1 _15311_/A sky130_fd_sc_hd__nor2_1
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16289_ _16533_/Q _16289_/D vssd1 vssd1 vccd1 vccd1 _16289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09801_ _09801_/A vssd1 vssd1 vccd1 vccd1 _10178_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07993_ _16615_/Q vssd1 vssd1 vccd1 vccd1 _14113_/A sky130_fd_sc_hd__inv_4
XFILLER_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09732_ _15685_/Q _09919_/B _09739_/C vssd1 vssd1 vccd1 vccd1 _09734_/B sky130_fd_sc_hd__and3_1
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09663_ _09663_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _15668_/D sky130_fd_sc_hd__nor2_1
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08614_ _13521_/A vssd1 vssd1 vccd1 vccd1 _10501_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ _09587_/C _09588_/C _09591_/Y _09598_/A vssd1 vssd1 vccd1 vccd1 _09598_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_82_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _08545_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _15315_/C sky130_fd_sc_hd__xor2_2
XFILLER_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08476_ _08476_/A _08492_/A vssd1 vssd1 vccd1 vccd1 _08477_/B sky130_fd_sc_hd__xor2_1
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09028_ _15542_/Q _09192_/B _09028_/C vssd1 vssd1 vccd1 vccd1 _09029_/B sky130_fd_sc_hd__and3_1
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13990_ _13990_/A _13997_/B vssd1 vssd1 vccd1 vccd1 _13992_/A sky130_fd_sc_hd__or2_1
XFILLER_19_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12941_ _12941_/A _12941_/B _12941_/C vssd1 vssd1 vccd1 vccd1 _12942_/C sky130_fd_sc_hd__nand3_1
XFILLER_58_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15660_ _15791_/CLK _15660_/D vssd1 vssd1 vccd1 vccd1 _15660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12872_ _12889_/C vssd1 vssd1 vccd1 vccd1 _12896_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14611_ _14895_/A vssd1 vssd1 vccd1 vccd1 _14839_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _11821_/Y _11817_/C _11819_/Y _11820_/X vssd1 vssd1 vccd1 vccd1 _11824_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _16570_/CLK _15591_/D vssd1 vssd1 vccd1 vccd1 _15591_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14540_/Y _14535_/C _14538_/Y _14549_/A vssd1 vssd1 vccd1 vccd1 _14549_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11754_/A vssd1 vssd1 vccd1 vccd1 _16015_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10809_/A _10705_/B _10709_/B vssd1 vssd1 vccd1 vccd1 _15863_/D sky130_fd_sc_hd__nor3_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _16402_/Q _14591_/B _14480_/C vssd1 vssd1 vccd1 vccd1 _14473_/Y sky130_fd_sc_hd__nand3_1
X_11685_ _11706_/C vssd1 vssd1 vccd1 vccd1 _11721_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16212_ _16237_/CLK _16212_/D vssd1 vssd1 vccd1 vccd1 _16212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13424_ _16253_/Q _13645_/B _13424_/C vssd1 vssd1 vccd1 vccd1 _13432_/B sky130_fd_sc_hd__and3_1
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10636_ _10649_/A _10636_/B _10636_/C vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__and3_1
XFILLER_127_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _16261_/CLK _16143_/D vssd1 vssd1 vccd1 vccd1 _16143_/Q sky130_fd_sc_hd__dfxtp_1
X_13355_ _13355_/A vssd1 vssd1 vccd1 vccd1 _16242_/D sky130_fd_sc_hd__clkbuf_1
X_10567_ _10567_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10569_/B sky130_fd_sc_hd__nor2_1
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ _12306_/A vssd1 vssd1 vccd1 vccd1 _16093_/D sky130_fd_sc_hd__clkbuf_1
X_16074_ _16118_/CLK _16074_/D vssd1 vssd1 vccd1 vccd1 _16074_/Q sky130_fd_sc_hd__dfxtp_1
X_13286_ _13302_/A _13286_/B _13286_/C vssd1 vssd1 vccd1 vccd1 _13287_/A sky130_fd_sc_hd__and3_1
X_10498_ _10498_/A vssd1 vssd1 vccd1 vccd1 _15825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15025_ _15025_/A vssd1 vssd1 vccd1 vccd1 _16489_/D sky130_fd_sc_hd__clkbuf_1
X_12237_ _12466_/A _12243_/C vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__or2_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12168_ _12165_/Y _12166_/X _12167_/Y _12163_/C vssd1 vssd1 vccd1 vccd1 _12170_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_123_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11119_ _11236_/A _11119_/B _11123_/A vssd1 vssd1 vccd1 vccd1 _15926_/D sky130_fd_sc_hd__nor3_1
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12099_ _16066_/Q _12210_/B _12100_/C vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__and3_1
X_15927_ _15365_/A _15927_/D vssd1 vssd1 vccd1 vccd1 _15927_/Q sky130_fd_sc_hd__dfxtp_1
Xinput6 io_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_4
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15858_ _16570_/CLK _15858_/D vssd1 vssd1 vccd1 vccd1 _15858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14809_ _14805_/Y _14807_/X _14808_/Y _14803_/C vssd1 vssd1 vccd1 vccd1 _14811_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_33_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15789_ _15791_/CLK _15789_/D vssd1 vssd1 vccd1 vccd1 _15789_/Q sky130_fd_sc_hd__dfxtp_1
X_08330_ _08330_/A _08330_/B vssd1 vssd1 vccd1 vccd1 _08336_/A sky130_fd_sc_hd__nand2_1
X_08261_ _15471_/Q vssd1 vssd1 vccd1 vccd1 _08590_/C sky130_fd_sc_hd__clkinv_2
XFILLER_20_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08192_ _10675_/C _07970_/B _08191_/X vssd1 vssd1 vccd1 vccd1 _08346_/B sky130_fd_sc_hd__o21a_2
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07976_ _15786_/Q vssd1 vssd1 vccd1 vccd1 _10178_/C sky130_fd_sc_hd__clkinv_4
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _15682_/Q _09739_/C _09714_/X vssd1 vssd1 vccd1 vccd1 _09718_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09646_ _09643_/A _09643_/B _09642_/Y _09645_/Y vssd1 vssd1 vccd1 vccd1 _15664_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09577_ _15669_/Q vssd1 vssd1 vccd1 vccd1 _09581_/C sky130_fd_sc_hd__inv_2
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08528_ _09126_/A vssd1 vssd1 vccd1 vccd1 _15312_/A sky130_fd_sc_hd__buf_2
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08459_ _08459_/A _08459_/B vssd1 vssd1 vccd1 vccd1 _08461_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11470_ _12886_/A vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__buf_4
XFILLER_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10421_ _15803_/Q _15802_/Q _15801_/Q _10227_/X vssd1 vssd1 vccd1 vccd1 _15813_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_136_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13140_ _13705_/A vssd1 vssd1 vccd1 vccd1 _13140_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10352_ _10399_/A _10352_/B _10352_/C vssd1 vssd1 vccd1 vccd1 _10353_/A sky130_fd_sc_hd__and3_1
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _13069_/Y _13065_/C _13067_/Y _13068_/X vssd1 vssd1 vccd1 vccd1 _13072_/C
+ sky130_fd_sc_hd__a211o_1
X_10283_ _10307_/B vssd1 vssd1 vccd1 vccd1 _10313_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_3_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12022_ _12038_/C vssd1 vssd1 vccd1 vccd1 _12045_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16761_ _16761_/A _07780_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
X_13973_ _16331_/Q _14193_/B _13981_/C vssd1 vssd1 vccd1 vccd1 _13973_/X sky130_fd_sc_hd__and3_1
XFILLER_101_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15712_ _15812_/CLK _15712_/D vssd1 vssd1 vccd1 vccd1 _15712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12924_ _12924_/A vssd1 vssd1 vccd1 vccd1 _13151_/A sky130_fd_sc_hd__clkbuf_2
X_16692_ _16692_/A _07790_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
X_15643_ _15791_/CLK _15643_/D vssd1 vssd1 vccd1 vccd1 _15643_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _12853_/Y _12847_/C _12851_/Y _12862_/A vssd1 vssd1 vccd1 vccd1 _12862_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _16024_/Q _11814_/C _11748_/X vssd1 vssd1 vccd1 vccd1 _11810_/B sky130_fd_sc_hd__a21o_1
X_15574_ _15812_/CLK _15574_/D vssd1 vssd1 vccd1 vccd1 _15574_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12783_/Y _12784_/X _12785_/Y _12781_/C vssd1 vssd1 vccd1 vccd1 _12788_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14521_/Y _14523_/X _14524_/Y _14519_/C vssd1 vssd1 vccd1 vccd1 _14527_/B
+ sky130_fd_sc_hd__o211ai_1
X_11737_ _11737_/A _11737_/B _11737_/C vssd1 vssd1 vccd1 vccd1 _11738_/C sky130_fd_sc_hd__or3_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14456_ _14456_/A vssd1 vssd1 vccd1 vccd1 _16399_/D sky130_fd_sc_hd__clkbuf_1
X_11668_ _16005_/Q _11668_/B _11668_/C vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__and3_1
X_13407_ _13407_/A vssd1 vssd1 vccd1 vccd1 _13631_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10619_ _10613_/B _10616_/B _10414_/X vssd1 vssd1 vccd1 vccd1 _10620_/B sky130_fd_sc_hd__o21a_1
X_14387_ _14669_/A vssd1 vssd1 vccd1 vccd1 _14387_/X sky130_fd_sc_hd__clkbuf_2
X_11599_ _15995_/Q _11607_/C _11485_/X vssd1 vssd1 vccd1 vccd1 _11599_/Y sky130_fd_sc_hd__a21oi_1
X_16126_ _16554_/Q _16126_/D vssd1 vssd1 vccd1 vccd1 _16126_/Q sky130_fd_sc_hd__dfxtp_2
X_13338_ _13332_/C _13333_/C _13335_/Y _13336_/X vssd1 vssd1 vccd1 vccd1 _13339_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16057_ _16118_/CLK _16057_/D vssd1 vssd1 vccd1 vccd1 _16057_/Q sky130_fd_sc_hd__dfxtp_1
X_13269_ _13269_/A vssd1 vssd1 vccd1 vccd1 _13283_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15008_ _15009_/B _15009_/C _14954_/X vssd1 vssd1 vccd1 vccd1 _15010_/B sky130_fd_sc_hd__o21ai_1
XFILLER_97_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07830_ _07830_/A vssd1 vssd1 vccd1 vccd1 _07830_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07761_ _07762_/A vssd1 vssd1 vccd1 vccd1 _07761_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09500_ _09501_/B _09501_/C _09501_/A vssd1 vssd1 vccd1 vccd1 _09502_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _09750_/A vssd1 vssd1 vccd1 vccd1 _09431_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ _10183_/A vssd1 vssd1 vccd1 vccd1 _09362_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_33_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ _08109_/C _08309_/Y _08312_/Y vssd1 vssd1 vccd1 vccd1 _15447_/D sky130_fd_sc_hd__o21a_1
X_09293_ _09698_/A vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_11 _08854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _07774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08244_ _08244_/A _08371_/A vssd1 vssd1 vccd1 vccd1 _08279_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_33 _14220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 _15415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08175_ _08176_/A _08176_/B vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07959_ _16609_/Q vssd1 vssd1 vccd1 vccd1 _13777_/A sky130_fd_sc_hd__inv_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10970_ _15905_/Q _11026_/B _10970_/C vssd1 vssd1 vccd1 vccd1 _10970_/Y sky130_fd_sc_hd__nand3_1
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09629_ _09629_/A vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__buf_2
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12640_ _12751_/A vssd1 vssd1 vccd1 vccd1 _12681_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12571_ _12568_/Y _12580_/A _12570_/Y _12565_/C vssd1 vssd1 vccd1 vccd1 _12573_/B
+ sky130_fd_sc_hd__o211a_1
X_14310_ _16379_/Q _14472_/B _14317_/C vssd1 vssd1 vccd1 vccd1 _14310_/X sky130_fd_sc_hd__and3_1
X_11522_ _12373_/A vssd1 vssd1 vccd1 vccd1 _11750_/B sky130_fd_sc_hd__clkbuf_2
X_15290_ _15291_/A _15291_/B vssd1 vssd1 vccd1 vccd1 _15292_/A sky130_fd_sc_hd__or2_1
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _14241_/A vssd1 vssd1 vccd1 vccd1 _16368_/D sky130_fd_sc_hd__clkbuf_1
X_11453_ _11491_/A _11453_/B _11453_/C vssd1 vssd1 vccd1 vccd1 _11454_/A sky130_fd_sc_hd__and3_1
X_10404_ _10401_/Y _10410_/A _10403_/Y _10399_/C vssd1 vssd1 vccd1 vccd1 _10406_/B
+ sky130_fd_sc_hd__o211a_1
X_14172_ _16360_/Q _14179_/C _14008_/X vssd1 vssd1 vccd1 vccd1 _14175_/B sky130_fd_sc_hd__a21o_1
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11384_ _11384_/A vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__clkbuf_2
X_13123_ _13131_/A _13123_/B _13123_/C vssd1 vssd1 vccd1 vccd1 _13124_/A sky130_fd_sc_hd__and3_1
X_10335_ _15799_/Q _10434_/B _10342_/C vssd1 vssd1 vccd1 vccd1 _10337_/C sky130_fd_sc_hd__nand3_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _13052_/Y _13053_/X _13049_/C _13050_/C vssd1 vssd1 vccd1 vccd1 _13056_/B
+ sky130_fd_sc_hd__o211ai_1
X_10266_ _15785_/Q _10267_/C _10104_/X vssd1 vssd1 vccd1 vccd1 _10268_/A sky130_fd_sc_hd__a21oi_1
XFILLER_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12005_ _12003_/Y _11998_/C _12001_/Y _12012_/A vssd1 vssd1 vccd1 vccd1 _12012_/B
+ sky130_fd_sc_hd__a211oi_1
X_10197_ _15774_/Q _10446_/B _10206_/C vssd1 vssd1 vccd1 vccd1 _10197_/X sky130_fd_sc_hd__and3_1
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16744_ _16744_/A _07760_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_13956_ _16329_/Q _13966_/C _13736_/X vssd1 vssd1 vccd1 vccd1 _13956_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12907_ _12907_/A _12907_/B _12907_/C vssd1 vssd1 vccd1 vccd1 _12908_/A sky130_fd_sc_hd__and3_1
X_13887_ _13900_/C vssd1 vssd1 vccd1 vccd1 _13908_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15626_ _15791_/CLK _15626_/D vssd1 vssd1 vccd1 vccd1 _15626_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _12836_/Y _12831_/C _12833_/Y _12835_/X vssd1 vssd1 vccd1 vccd1 _12839_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_62_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12769_ _16161_/Q _12778_/C _12605_/X vssd1 vssd1 vccd1 vccd1 _12769_/Y sky130_fd_sc_hd__a21oi_1
X_15557_ _16551_/CLK _15557_/D vssd1 vssd1 vccd1 vccd1 _15557_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14508_ _16409_/Q _14516_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14511_/B sky130_fd_sc_hd__a21o_1
X_15488_ _16570_/CLK _15488_/D vssd1 vssd1 vccd1 vccd1 _15488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14439_ _14439_/A vssd1 vssd1 vccd1 vccd1 _14476_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16109_ _16554_/Q _16109_/D vssd1 vssd1 vccd1 vccd1 _16109_/Q sky130_fd_sc_hd__dfxtp_1
X_09980_ _09980_/A _09980_/B vssd1 vssd1 vccd1 vccd1 _15731_/D sky130_fd_sc_hd__nor2_1
X_08931_ _15534_/Q vssd1 vssd1 vccd1 vccd1 _08937_/C sky130_fd_sc_hd__inv_2
XFILLER_130_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08862_ _08860_/Y _08868_/A _08851_/C _08852_/C vssd1 vssd1 vccd1 vccd1 _08864_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07813_ _07837_/A vssd1 vssd1 vccd1 vccd1 _07818_/A sky130_fd_sc_hd__buf_12
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08793_ _08793_/A _08793_/B vssd1 vssd1 vccd1 vccd1 _15487_/D sky130_fd_sc_hd__nor2_1
XFILLER_123_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09414_ _09414_/A vssd1 vssd1 vccd1 vccd1 _15617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09345_ _09339_/Y _09340_/X _09342_/B vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__o21a_1
XFILLER_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09276_ _09276_/A _09276_/B vssd1 vssd1 vccd1 vccd1 _09276_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08227_ _08227_/A _08348_/A vssd1 vssd1 vccd1 vccd1 _08283_/A sky130_fd_sc_hd__xnor2_4
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08158_ _08353_/A _08158_/B vssd1 vssd1 vccd1 vccd1 _08330_/B sky130_fd_sc_hd__and2_1
XFILLER_107_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08089_ _16592_/Q _08270_/B vssd1 vssd1 vccd1 vccd1 _08090_/B sky130_fd_sc_hd__xnor2_1
XFILLER_122_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ _10124_/C vssd1 vssd1 vccd1 vccd1 _10133_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10051_ _15748_/Q _10307_/C _10051_/C vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__and3_1
XFILLER_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13810_ _13808_/Y _13803_/C _13805_/Y _13806_/X vssd1 vssd1 vccd1 vccd1 _13811_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14790_ _16453_/Q _14790_/B _14800_/C vssd1 vssd1 vccd1 vccd1 _14795_/A sky130_fd_sc_hd__and3_1
XFILLER_91_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13741_ _13756_/A _13741_/B _13741_/C vssd1 vssd1 vccd1 vccd1 _13742_/A sky130_fd_sc_hd__and3_1
X_10953_ _15903_/Q _11118_/B _10963_/C vssd1 vssd1 vccd1 vccd1 _10959_/A sky130_fd_sc_hd__and3_1
XFILLER_73_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13672_ _13672_/A vssd1 vssd1 vccd1 vccd1 _16287_/D sky130_fd_sc_hd__clkbuf_1
X_16460_ input11/X _16460_/D vssd1 vssd1 vccd1 vccd1 _16460_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10884_ _11051_/A vssd1 vssd1 vccd1 vccd1 _10925_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15411_ _16165_/Q _16164_/Q _16163_/Q _15409_/X vssd1 vssd1 vccd1 vccd1 _16591_/D
+ sky130_fd_sc_hd__o31a_1
X_12623_ _12620_/Y _12621_/X _12622_/Y _12617_/C vssd1 vssd1 vccd1 vccd1 _12625_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16391_ input11/X _16391_/D vssd1 vssd1 vccd1 vccd1 _16391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15342_ _15340_/Y _15348_/A _15337_/C _15338_/C vssd1 vssd1 vccd1 vccd1 _15344_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12554_ _16129_/Q _12726_/B _12554_/C vssd1 vssd1 vccd1 vccd1 _12554_/Y sky130_fd_sc_hd__nand3_1
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11505_ _11503_/A _11503_/B _11504_/X vssd1 vssd1 vccd1 vccd1 _15980_/D sky130_fd_sc_hd__a21oi_1
X_15273_ _15274_/B _15274_/C _09207_/A vssd1 vssd1 vccd1 vccd1 _15275_/B sky130_fd_sc_hd__o21ai_1
X_12485_ _12485_/A vssd1 vssd1 vccd1 vccd1 _16119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14224_ _14245_/C vssd1 vssd1 vccd1 vccd1 _14260_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11436_ _15972_/Q _11607_/B _11436_/C vssd1 vssd1 vccd1 vccd1 _11446_/A sky130_fd_sc_hd__and3_1
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14155_ _14155_/A _14162_/B vssd1 vssd1 vccd1 vccd1 _14157_/A sky130_fd_sc_hd__or2_1
X_11367_ _15963_/Q _11367_/B _11375_/C vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__and3_1
XFILLER_98_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13106_ _13107_/B _13107_/C _13107_/A vssd1 vssd1 vccd1 vccd1 _13108_/B sky130_fd_sc_hd__a21o_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _10318_/A _10318_/B vssd1 vssd1 vccd1 vccd1 _10319_/B sky130_fd_sc_hd__nor2_1
X_14086_ _14647_/A vssd1 vssd1 vccd1 vccd1 _14311_/B sky130_fd_sc_hd__clkbuf_2
X_11298_ _11319_/A _11298_/B _11298_/C vssd1 vssd1 vccd1 vccd1 _11299_/A sky130_fd_sc_hd__and3_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _13072_/A _13037_/B _13037_/C vssd1 vssd1 vccd1 vccd1 _13038_/A sky130_fd_sc_hd__and3_1
X_10249_ _10240_/C _10241_/C _10244_/Y _10247_/X vssd1 vssd1 vccd1 vccd1 _10250_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14988_ _16484_/Q _15041_/B _14995_/C vssd1 vssd1 vccd1 vccd1 _14988_/X sky130_fd_sc_hd__and3_1
XFILLER_75_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16727_ _16727_/A _07832_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13939_ _13997_/A _13939_/B _13939_/C vssd1 vssd1 vccd1 vccd1 _13940_/C sky130_fd_sc_hd__or3_1
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _15812_/CLK _15609_/D vssd1 vssd1 vccd1 vccd1 _15609_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16589_ _16595_/CLK _16589_/D vssd1 vssd1 vccd1 vccd1 _16589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09130_ _09006_/X _09128_/A _09129_/X vssd1 vssd1 vccd1 vccd1 _09130_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09061_ _09061_/A vssd1 vssd1 vccd1 vccd1 _15545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08012_ _16559_/Q _08218_/A _08012_/C vssd1 vssd1 vccd1 vccd1 _08218_/B sky130_fd_sc_hd__nand3_1
XFILLER_144_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09963_ _09962_/X _09961_/Y _08700_/A vssd1 vssd1 vccd1 vccd1 _09963_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08914_ _09117_/A vssd1 vssd1 vccd1 vccd1 _08914_/X sky130_fd_sc_hd__buf_2
XFILLER_131_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _10716_/A vssd1 vssd1 vccd1 vccd1 _09894_/X sky130_fd_sc_hd__buf_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08845_ _15503_/Q _08845_/B _08849_/C vssd1 vssd1 vccd1 vccd1 _08851_/A sky130_fd_sc_hd__and3_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08776_ _08846_/A _08776_/B _08781_/B vssd1 vssd1 vccd1 vccd1 _15483_/D sky130_fd_sc_hd__nor3_1
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09328_ _15603_/Q _09329_/C _15341_/B vssd1 vssd1 vccd1 vccd1 _09328_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ _15593_/Q _09364_/B _09267_/C vssd1 vssd1 vccd1 vccd1 _09261_/C sky130_fd_sc_hd__nand3_1
XFILLER_127_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _16090_/Q _12493_/B _12271_/C vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__and3_1
XFILLER_107_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11221_ _11332_/A _11226_/C vssd1 vssd1 vccd1 vccd1 _11221_/X sky130_fd_sc_hd__or2_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11152_ _15932_/Q _11322_/B _11152_/C vssd1 vssd1 vccd1 vccd1 _11163_/A sky130_fd_sc_hd__and3_1
X_10103_ _10179_/A _10103_/B _10108_/B vssd1 vssd1 vccd1 vccd1 _15755_/D sky130_fd_sc_hd__nor3_1
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15960_ _16005_/CLK _15960_/D vssd1 vssd1 vccd1 vccd1 _15960_/Q sky130_fd_sc_hd__dfxtp_1
X_11083_ _15923_/Q _11093_/C _10919_/X vssd1 vssd1 vccd1 vccd1 _11083_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10034_ _10034_/A _10034_/B _10034_/C vssd1 vssd1 vccd1 vccd1 _10035_/C sky130_fd_sc_hd__nand3_1
X_14911_ _14911_/A vssd1 vssd1 vccd1 vccd1 _15129_/B sky130_fd_sc_hd__buf_2
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15891_ _16553_/Q _15891_/D vssd1 vssd1 vccd1 vccd1 _15891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14842_ _16397_/Q _16396_/Q _16395_/Q _14615_/X vssd1 vssd1 vccd1 vccd1 _16460_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_64_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14773_ _15058_/A vssd1 vssd1 vccd1 vccd1 _15005_/A sky130_fd_sc_hd__clkbuf_2
X_11985_ _12269_/A vssd1 vssd1 vccd1 vccd1 _12210_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16512_ _16607_/CLK _16512_/D vssd1 vssd1 vccd1 vccd1 _16512_/Q sky130_fd_sc_hd__dfxtp_1
X_13724_ _16295_/Q _13765_/C _13495_/X vssd1 vssd1 vccd1 vccd1 _13727_/B sky130_fd_sc_hd__a21oi_1
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10936_ _10936_/A _10936_/B vssd1 vssd1 vccd1 vccd1 _10937_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16443_ _16607_/CLK _16443_/D vssd1 vssd1 vccd1 vccd1 _16443_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10867_ _15892_/Q _10878_/C _10866_/X vssd1 vssd1 vccd1 vccd1 _10867_/Y sky130_fd_sc_hd__a21oi_1
X_13655_ _13656_/B _13656_/C _13546_/X vssd1 vssd1 vccd1 vccd1 _13657_/B sky130_fd_sc_hd__o21ai_1
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _16137_/Q _12614_/C _12605_/X vssd1 vssd1 vccd1 vccd1 _12606_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16374_ _16389_/CLK _16374_/D vssd1 vssd1 vccd1 vccd1 _16374_/Q sky130_fd_sc_hd__dfxtp_2
X_13586_ _16276_/Q _13586_/B _13586_/C vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__and3_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _15881_/Q _10922_/B _10805_/C vssd1 vssd1 vccd1 vccd1 _10798_/Y sky130_fd_sc_hd__nand3_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15325_ _15324_/Y _15312_/B _15316_/B _15322_/Y _15320_/Y vssd1 vssd1 vccd1 vccd1
+ _15325_/X sky130_fd_sc_hd__a311o_1
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12537_ _16128_/Q _12545_/C _12316_/X vssd1 vssd1 vccd1 vccd1 _12540_/B sky130_fd_sc_hd__a21o_1
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15256_ _15253_/Y _15254_/X _15255_/Y _15251_/C vssd1 vssd1 vccd1 vccd1 _15258_/B
+ sky130_fd_sc_hd__o211ai_1
X_12468_ _12468_/A vssd1 vssd1 vccd1 vccd1 _12505_/A sky130_fd_sc_hd__clkbuf_2
X_11419_ _15970_/Q _11644_/B _11420_/C vssd1 vssd1 vccd1 vccd1 _11419_/X sky130_fd_sc_hd__and3_1
X_14207_ _16365_/Q _14207_/B _14207_/C vssd1 vssd1 vccd1 vccd1 _14217_/B sky130_fd_sc_hd__and3_1
X_15187_ _16518_/Q _15195_/C _10782_/B vssd1 vssd1 vccd1 vccd1 _15187_/Y sky130_fd_sc_hd__a21oi_1
X_12399_ _12399_/A vssd1 vssd1 vccd1 vccd1 _16106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14138_ _14145_/A _14138_/B _14138_/C vssd1 vssd1 vccd1 vccd1 _14139_/A sky130_fd_sc_hd__and3_1
XFILLER_99_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14069_ _14090_/A _14069_/B _14069_/C vssd1 vssd1 vccd1 vccd1 _14070_/A sky130_fd_sc_hd__and3_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ _09076_/A vssd1 vssd1 vccd1 vccd1 _08630_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08561_ _15453_/Q _08561_/B vssd1 vssd1 vccd1 vccd1 _08568_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08492_ _08492_/A _08476_/A vssd1 vssd1 vccd1 vccd1 _08492_/X sky130_fd_sc_hd__or2b_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09113_ _10060_/A vssd1 vssd1 vccd1 vccd1 _09849_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09044_ _09044_/A _09044_/B vssd1 vssd1 vccd1 vccd1 _15541_/D sky130_fd_sc_hd__nor2_1
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09946_ _09946_/A _09946_/B _09950_/A vssd1 vssd1 vccd1 vccd1 _15724_/D sky130_fd_sc_hd__nor3_1
XFILLER_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _15712_/Q _09884_/C _09683_/X vssd1 vssd1 vccd1 vccd1 _09880_/A sky130_fd_sc_hd__a21oi_1
XFILLER_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08828_ _08823_/B _08826_/B _08698_/X vssd1 vssd1 vccd1 vccd1 _08836_/C sky130_fd_sc_hd__o21a_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _08766_/C vssd1 vssd1 vccd1 vccd1 _08779_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _12901_/A vssd1 vssd1 vccd1 vccd1 _11770_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _15885_/Q vssd1 vssd1 vccd1 vccd1 _10726_/C sky130_fd_sc_hd__inv_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13440_ _13725_/A vssd1 vssd1 vccd1 vccd1 _13665_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10652_ _15856_/Q _10652_/B _10652_/C vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__and3_1
XFILLER_41_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13371_ _13371_/A vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10583_ _15843_/Q _10726_/B _10583_/C vssd1 vssd1 vccd1 vccd1 _10588_/A sky130_fd_sc_hd__and3_1
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15110_ _15110_/A _15117_/B vssd1 vssd1 vccd1 vccd1 _15112_/A sky130_fd_sc_hd__or2_1
X_12322_ _12322_/A vssd1 vssd1 vccd1 vccd1 _16095_/D sky130_fd_sc_hd__clkbuf_1
X_16090_ _16118_/CLK _16090_/D vssd1 vssd1 vccd1 vccd1 _16090_/Q sky130_fd_sc_hd__dfxtp_1
X_15041_ _16493_/Q _15041_/B _15049_/C vssd1 vssd1 vccd1 vccd1 _15041_/X sky130_fd_sc_hd__and3_1
XFILLER_107_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12253_ _12371_/A _12253_/B _12257_/A vssd1 vssd1 vccd1 vccd1 _16086_/D sky130_fd_sc_hd__nor3_1
XFILLER_108_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11204_ _15939_/Q _11367_/B _11211_/C vssd1 vssd1 vccd1 vccd1 _11204_/X sky130_fd_sc_hd__and3_1
XFILLER_123_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ _12182_/A _12182_/B _12183_/X vssd1 vssd1 vccd1 vccd1 _16076_/D sky130_fd_sc_hd__a21oi_1
XFILLER_123_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11135_ _12269_/A vssd1 vssd1 vccd1 vccd1 _11359_/B sky130_fd_sc_hd__buf_2
XFILLER_110_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15943_ _15365_/A _15943_/D vssd1 vssd1 vccd1 vccd1 _15943_/Q sky130_fd_sc_hd__dfxtp_1
X_11066_ _11066_/A _11066_/B _11066_/C vssd1 vssd1 vccd1 vccd1 _11067_/C sky130_fd_sc_hd__nand3_1
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10017_ _10017_/A _10017_/B vssd1 vssd1 vccd1 vccd1 _10017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15874_ _16570_/CLK _15874_/D vssd1 vssd1 vccd1 vccd1 _15874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14825_ _14822_/Y _14833_/A _14824_/Y _14819_/C vssd1 vssd1 vccd1 vccd1 _14827_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14756_ _16448_/Q _14756_/B _14764_/C vssd1 vssd1 vccd1 vccd1 _14756_/X sky130_fd_sc_hd__and3_1
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11968_ _16047_/Q _12010_/C _11802_/X vssd1 vssd1 vccd1 vccd1 _11970_/B sky130_fd_sc_hd__a21oi_1
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13707_ input6/X vssd1 vssd1 vccd1 vccd1 _14830_/A sky130_fd_sc_hd__buf_4
X_10919_ _12968_/A vssd1 vssd1 vccd1 vccd1 _10919_/X sky130_fd_sc_hd__buf_2
X_11899_ _11899_/A _11899_/B vssd1 vssd1 vccd1 vccd1 _11900_/B sky130_fd_sc_hd__nor2_1
X_14687_ _14687_/A vssd1 vssd1 vccd1 vccd1 _16435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16426_ _16595_/CLK _16426_/D vssd1 vssd1 vccd1 vccd1 _16426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ _13638_/A vssd1 vssd1 vccd1 vccd1 _13869_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16357_ _16389_/CLK _16357_/D vssd1 vssd1 vccd1 vccd1 _16357_/Q sky130_fd_sc_hd__dfxtp_1
X_13569_ _13569_/A vssd1 vssd1 vccd1 vccd1 _16272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ _16709_/A _15321_/B _15307_/C vssd1 vssd1 vccd1 vccd1 _15309_/B sky130_fd_sc_hd__a21oi_1
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16288_ _16533_/Q _16288_/D vssd1 vssd1 vccd1 vccd1 _16288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15239_ _15239_/A vssd1 vssd1 vccd1 vccd1 _16525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09800_ _15699_/Q _09845_/C _09714_/X vssd1 vssd1 vccd1 vccd1 _09803_/B sky130_fd_sc_hd__a21oi_1
XFILLER_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07992_ _07992_/A _08204_/B vssd1 vssd1 vccd1 vccd1 _08208_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09731_ _15685_/Q _09739_/C _09683_/X vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__a21oi_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09662_ _09617_/X _09486_/X _09656_/B _09487_/X vssd1 vssd1 vccd1 vccd1 _09663_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08613_ _13288_/A vssd1 vssd1 vccd1 vccd1 _13521_/A sky130_fd_sc_hd__buf_8
X_09593_ _09591_/Y _09598_/A _09587_/C _09588_/C vssd1 vssd1 vccd1 vccd1 _09595_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _08556_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__xor2_2
XFILLER_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08475_ _08475_/A _08475_/B vssd1 vssd1 vccd1 vccd1 _08492_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09027_ _10501_/A vssd1 vssd1 vccd1 vccd1 _09192_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_123_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09929_ _09924_/Y _09927_/X _09928_/Y vssd1 vssd1 vccd1 vccd1 _15719_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12940_ _12941_/B _12941_/C _12941_/A vssd1 vssd1 vccd1 vccd1 _12942_/B sky130_fd_sc_hd__a21o_1
XFILLER_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12871_ _16593_/Q vssd1 vssd1 vccd1 vccd1 _12889_/C sky130_fd_sc_hd__inv_2
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14610_ _14612_/B _14612_/C _14387_/X vssd1 vssd1 vccd1 vccd1 _14613_/B sky130_fd_sc_hd__o21ai_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11819_/Y _11820_/X _11821_/Y _11817_/C vssd1 vssd1 vccd1 vccd1 _11824_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15590_ _16570_/CLK _15590_/D vssd1 vssd1 vccd1 vccd1 _15590_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _11776_/A _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11754_/A sky130_fd_sc_hd__and3_1
X_14541_ _14538_/Y _14549_/A _14540_/Y _14535_/C vssd1 vssd1 vccd1 vccd1 _14543_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10702_/Y _10695_/C _10699_/Y _10709_/A vssd1 vssd1 vccd1 vccd1 _10709_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11684_ _11698_/C vssd1 vssd1 vccd1 vccd1 _11706_/C sky130_fd_sc_hd__clkbuf_1
X_14472_ _16403_/Q _14472_/B _14480_/C vssd1 vssd1 vccd1 vccd1 _14472_/X sky130_fd_sc_hd__and3_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _16237_/CLK _16211_/D vssd1 vssd1 vccd1 vccd1 _16211_/Q sky130_fd_sc_hd__dfxtp_1
X_10635_ _10635_/A _10635_/B _10635_/C vssd1 vssd1 vccd1 vccd1 _10636_/C sky130_fd_sc_hd__nand3_1
X_13423_ _13423_/A vssd1 vssd1 vccd1 vccd1 _13645_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16142_ _16261_/CLK _16142_/D vssd1 vssd1 vccd1 vccd1 _16142_/Q sky130_fd_sc_hd__dfxtp_2
X_13354_ _13354_/A _13354_/B _13354_/C vssd1 vssd1 vccd1 vccd1 _13355_/A sky130_fd_sc_hd__and3_1
XFILLER_6_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10566_ _10566_/A _10566_/B vssd1 vssd1 vccd1 vccd1 _10569_/A sky130_fd_sc_hd__or2_1
XFILLER_139_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12305_ _12343_/A _12305_/B _12305_/C vssd1 vssd1 vccd1 vccd1 _12306_/A sky130_fd_sc_hd__and3_1
XFILLER_6_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13285_ _13279_/C _13280_/C _13282_/Y _13283_/X vssd1 vssd1 vccd1 vccd1 _13286_/C
+ sky130_fd_sc_hd__a211o_1
X_16073_ _16118_/CLK _16073_/D vssd1 vssd1 vccd1 vccd1 _16073_/Q sky130_fd_sc_hd__dfxtp_1
X_10497_ _10497_/A _10497_/B _10497_/C vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__and3_1
XFILLER_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _12236_/A _12236_/B vssd1 vssd1 vccd1 vccd1 _12243_/C sky130_fd_sc_hd__nor2_1
X_15024_ _15045_/A _15024_/B _15024_/C vssd1 vssd1 vccd1 vccd1 _15025_/A sky130_fd_sc_hd__and3_1
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12167_ _16074_/Q _12340_/B _12173_/C vssd1 vssd1 vccd1 vccd1 _12167_/Y sky130_fd_sc_hd__nand3_1
XFILLER_111_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11118_ _15927_/Q _11118_/B _11128_/C vssd1 vssd1 vccd1 vccd1 _11123_/A sky130_fd_sc_hd__and3_1
XFILLER_49_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12098_ _16066_/Q _12100_/C _11875_/X vssd1 vssd1 vccd1 vccd1 _12098_/Y sky130_fd_sc_hd__a21oi_1
X_16685__90 vssd1 vssd1 vccd1 vccd1 _16685__90/HI _16761_/A sky130_fd_sc_hd__conb_1
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15926_ _15365_/A _15926_/D vssd1 vssd1 vccd1 vccd1 _15926_/Q sky130_fd_sc_hd__dfxtp_2
X_11049_ _11049_/A _11053_/C vssd1 vssd1 vccd1 vccd1 _11049_/X sky130_fd_sc_hd__or2_1
Xinput7 io_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XFILLER_37_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15857_ _16570_/CLK _15857_/D vssd1 vssd1 vccd1 vccd1 _15857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _16455_/Q _14982_/B _14808_/C vssd1 vssd1 vccd1 vccd1 _14808_/Y sky130_fd_sc_hd__nand3_1
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15788_ _15791_/CLK _15788_/D vssd1 vssd1 vccd1 vccd1 _15788_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14739_ _14760_/A _14739_/B _14739_/C vssd1 vssd1 vccd1 vccd1 _14740_/A sky130_fd_sc_hd__and3_1
XFILLER_60_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ _08458_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08386_/A sky130_fd_sc_hd__nand2_2
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16409_ input11/X _16409_/D vssd1 vssd1 vccd1 vccd1 _16409_/Q sky130_fd_sc_hd__dfxtp_1
X_08191_ _10767_/A _08191_/B vssd1 vssd1 vccd1 vccd1 _08191_/X sky130_fd_sc_hd__or2_1
XFILLER_9_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07975_ _15768_/Q vssd1 vssd1 vccd1 vccd1 _10076_/C sky130_fd_sc_hd__clkinv_4
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _09943_/A vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _09643_/X _09642_/Y _09644_/X vssd1 vssd1 vccd1 vccd1 _09645_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09576_ _15641_/Q _15640_/Q _15639_/Q _09536_/X vssd1 vssd1 vccd1 vccd1 _15651_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _10430_/A vssd1 vssd1 vccd1 vccd1 _09126_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ _08458_/A _08458_/B vssd1 vssd1 vccd1 vccd1 _08459_/B sky130_fd_sc_hd__or2_1
XFILLER_50_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08389_ _08268_/A _08268_/B _08459_/A _08388_/X vssd1 vssd1 vccd1 vccd1 _08458_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_137_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10420_ _10276_/X _10416_/B _10419_/Y vssd1 vssd1 vccd1 vccd1 _15812_/D sky130_fd_sc_hd__o21a_1
XFILLER_137_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10351_ _10349_/Y _10345_/C _10347_/Y _10348_/X vssd1 vssd1 vccd1 vccd1 _10352_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_3_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13070_ _13067_/Y _13068_/X _13069_/Y _13065_/C vssd1 vssd1 vccd1 vccd1 _13072_/B
+ sky130_fd_sc_hd__o211ai_1
X_10282_ _10294_/B vssd1 vssd1 vccd1 vccd1 _10307_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12021_ _16578_/Q vssd1 vssd1 vccd1 vccd1 _12038_/C sky130_fd_sc_hd__inv_2
XFILLER_105_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16760_ _16760_/A _07779_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
X_13972_ _14814_/A vssd1 vssd1 vccd1 vccd1 _14193_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15711_ _15812_/CLK _15711_/D vssd1 vssd1 vccd1 vccd1 _15711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12923_ _12925_/B _12925_/C _12699_/X vssd1 vssd1 vccd1 vccd1 _12926_/B sky130_fd_sc_hd__o21ai_1
X_16691_ _16691_/A _07789_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_46_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15642_ _15812_/CLK _15642_/D vssd1 vssd1 vccd1 vccd1 _15642_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _12851_/Y _12862_/A _12853_/Y _12847_/C vssd1 vssd1 vccd1 vccd1 _12856_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _11805_/A _11805_/B _11810_/A vssd1 vssd1 vccd1 vccd1 _16022_/D sky130_fd_sc_hd__nor3_1
XFILLER_92_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15573_ _15812_/CLK _15573_/D vssd1 vssd1 vccd1 vccd1 _15573_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _16162_/Q _12904_/B _12792_/C vssd1 vssd1 vccd1 vccd1 _12785_/Y sky130_fd_sc_hd__nand3_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _16410_/Q _14697_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _14524_/Y sky130_fd_sc_hd__nand3_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11736_ _11737_/B _11737_/C _11567_/X vssd1 vssd1 vccd1 vccd1 _11738_/B sky130_fd_sc_hd__o21ai_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14455_ _14476_/A _14455_/B _14455_/C vssd1 vssd1 vccd1 vccd1 _14456_/A sky130_fd_sc_hd__and3_1
X_11667_ _16005_/Q _11668_/C _11441_/X vssd1 vssd1 vccd1 vccd1 _11669_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13406_ _16251_/Q _13416_/C _13184_/X vssd1 vssd1 vccd1 vccd1 _13406_/Y sky130_fd_sc_hd__a21oi_1
X_10618_ _10618_/A vssd1 vssd1 vccd1 vccd1 _15353_/A sky130_fd_sc_hd__buf_2
X_11598_ _11598_/A vssd1 vssd1 vccd1 vccd1 _15993_/D sky130_fd_sc_hd__clkbuf_1
X_14386_ _14439_/A vssd1 vssd1 vccd1 vccd1 _14424_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16125_ _16554_/Q _16125_/D vssd1 vssd1 vccd1 vccd1 _16125_/Q sky130_fd_sc_hd__dfxtp_1
X_13337_ _13335_/Y _13336_/X _13332_/C _13333_/C vssd1 vssd1 vccd1 vccd1 _13339_/B
+ sky130_fd_sc_hd__o211ai_1
X_10549_ _10589_/A _10549_/B _10549_/C vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__and3_1
XFILLER_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16056_ _16118_/CLK _16056_/D vssd1 vssd1 vccd1 vccd1 _16056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13268_ _13268_/A vssd1 vssd1 vccd1 vccd1 _16229_/D sky130_fd_sc_hd__clkbuf_1
X_15007_ _15007_/A vssd1 vssd1 vccd1 vccd1 _15045_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12219_ _16082_/Q _12340_/B _12226_/C vssd1 vssd1 vccd1 vccd1 _12219_/Y sky130_fd_sc_hd__nand3_1
X_13199_ _16221_/Q _13364_/B _13199_/C vssd1 vssd1 vccd1 vccd1 _13209_/B sky130_fd_sc_hd__and3_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07760_ _07762_/A vssd1 vssd1 vccd1 vccd1 _07760_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15909_ _15365_/A _15909_/D vssd1 vssd1 vccd1 vccd1 _15909_/Q sky130_fd_sc_hd__dfxtp_1
X_09430_ _09428_/X _09430_/B vssd1 vssd1 vccd1 vccd1 _09430_/X sky130_fd_sc_hd__and2b_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _09374_/A _09361_/B _09366_/A vssd1 vssd1 vccd1 vccd1 _15607_/D sky130_fd_sc_hd__nor3_1
XFILLER_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08312_ _08109_/C _08309_/Y _15344_/A vssd1 vssd1 vccd1 vccd1 _08312_/Y sky130_fd_sc_hd__a21oi_1
X_09292_ _09282_/Y _09286_/X _09288_/B vssd1 vssd1 vccd1 vccd1 _09295_/B sky130_fd_sc_hd__o21a_1
XANTENNA_12 _10393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _10755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08243_/A _08370_/A vssd1 vssd1 vccd1 vccd1 _08371_/A sky130_fd_sc_hd__xor2_4
XFILLER_138_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_34 _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08174_ _08328_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08176_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07958_ _12646_/A _07958_/B vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__xnor2_4
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07889_ _13097_/A _07889_/B vssd1 vssd1 vccd1 vccd1 _08132_/B sky130_fd_sc_hd__xnor2_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09628_ _15665_/Q _09636_/C _09583_/X vssd1 vssd1 vccd1 vccd1 _09632_/B sky130_fd_sc_hd__a21o_1
XFILLER_55_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09559_ _09557_/A _09557_/B _09556_/Y _09558_/Y vssd1 vssd1 vccd1 vccd1 _15646_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12570_ _16131_/Q _12629_/B _12578_/C vssd1 vssd1 vccd1 vccd1 _12570_/Y sky130_fd_sc_hd__nand3_1
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ _15984_/Q _11529_/C _11463_/X vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__a21o_1
XFILLER_11_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11452_ _11452_/A _11452_/B _11452_/C vssd1 vssd1 vccd1 vccd1 _11453_/C sky130_fd_sc_hd__or3_1
X_14240_ _14256_/A _14240_/B _14240_/C vssd1 vssd1 vccd1 vccd1 _14241_/A sky130_fd_sc_hd__and3_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10403_ _15810_/Q _10458_/B _10408_/C vssd1 vssd1 vccd1 vccd1 _10403_/Y sky130_fd_sc_hd__nand3_1
X_14171_ _14205_/A _14171_/B _14175_/A vssd1 vssd1 vccd1 vccd1 _16358_/D sky130_fd_sc_hd__nor3_1
X_11383_ _11383_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__nor2_1
X_10334_ _15799_/Q _10342_/C _10181_/X vssd1 vssd1 vccd1 vccd1 _10337_/B sky130_fd_sc_hd__a21o_1
X_13122_ _13120_/Y _13115_/C _13117_/Y _13119_/X vssd1 vssd1 vccd1 vccd1 _13123_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13053_ _16201_/Q _13053_/B _13053_/C vssd1 vssd1 vccd1 vccd1 _13053_/X sky130_fd_sc_hd__and3_1
XFILLER_127_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10265_ _10311_/A _10265_/B _10269_/B vssd1 vssd1 vccd1 vccd1 _15782_/D sky130_fd_sc_hd__nor3_1
XFILLER_87_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12004_ _12001_/Y _12012_/A _12003_/Y _11998_/C vssd1 vssd1 vccd1 vccd1 _12006_/B
+ sky130_fd_sc_hd__o211a_1
X_10196_ _10501_/A vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_120_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16655__60 vssd1 vssd1 vccd1 vccd1 _16655__60/HI _16731_/A sky130_fd_sc_hd__conb_1
XFILLER_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16743_ _16743_/A _07759_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_13955_ _13955_/A vssd1 vssd1 vccd1 vccd1 _16327_/D sky130_fd_sc_hd__clkbuf_1
X_12906_ _12904_/Y _12899_/C _12902_/Y _12903_/X vssd1 vssd1 vccd1 vccd1 _12907_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_62_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _13886_/A vssd1 vssd1 vccd1 vccd1 _13900_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15625_ _15791_/CLK _15625_/D vssd1 vssd1 vccd1 vccd1 _15625_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12833_/Y _12835_/X _12836_/Y _12831_/C vssd1 vssd1 vccd1 vccd1 _12839_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_22_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _15791_/CLK _15556_/D vssd1 vssd1 vccd1 vccd1 _15556_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12768_/A vssd1 vssd1 vccd1 vccd1 _16159_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14624_/A _14507_/B _14511_/A vssd1 vssd1 vccd1 vccd1 _16407_/D sky130_fd_sc_hd__nor3_1
X_11719_ _12567_/A vssd1 vssd1 vccd1 vccd1 _11719_/X sky130_fd_sc_hd__clkbuf_2
X_15487_ _16570_/CLK _15487_/D vssd1 vssd1 vccd1 vccd1 _15487_/Q sky130_fd_sc_hd__dfxtp_1
X_12699_ _13264_/A vssd1 vssd1 vccd1 vccd1 _12699_/X sky130_fd_sc_hd__clkbuf_2
Xinput10 io_in[9] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_4
X_14438_ _14436_/A _14436_/B _14437_/X vssd1 vssd1 vccd1 vccd1 _16396_/D sky130_fd_sc_hd__a21oi_1
XFILLER_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14369_ _14369_/A _14369_/B _14369_/C vssd1 vssd1 vccd1 vccd1 _14370_/A sky130_fd_sc_hd__and3_1
XFILLER_143_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16108_ _16554_/Q _16108_/D vssd1 vssd1 vccd1 vccd1 _16108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08930_ _15506_/Q _15505_/Q _15504_/Q _08887_/X vssd1 vssd1 vccd1 vccd1 _15516_/D
+ sky130_fd_sc_hd__o31a_1
X_16039_ _16118_/CLK _16039_/D vssd1 vssd1 vccd1 vccd1 _16039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08861_ _15505_/Q _08943_/B _08866_/C vssd1 vssd1 vccd1 vccd1 _08868_/A sky130_fd_sc_hd__and3_1
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07812_ input1/X vssd1 vssd1 vccd1 vccd1 _07837_/A sky130_fd_sc_hd__buf_4
X_08792_ _08706_/X _08790_/A _08708_/X vssd1 vssd1 vccd1 vccd1 _08793_/B sky130_fd_sc_hd__o21ai_1
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _09588_/A _09413_/B _09413_/C vssd1 vssd1 vccd1 vccd1 _09414_/A sky130_fd_sc_hd__and3_1
X_09344_ _09339_/Y _09342_/X _09343_/Y vssd1 vssd1 vccd1 vccd1 _15602_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ _15595_/Q _09837_/A _09286_/C vssd1 vssd1 vccd1 vccd1 _09277_/B sky130_fd_sc_hd__and3_1
XFILLER_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08226_ _08226_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _08348_/A sky130_fd_sc_hd__xnor2_2
X_08157_ _08157_/A _08157_/B vssd1 vssd1 vccd1 vccd1 _08158_/B sky130_fd_sc_hd__or2_1
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08088_ _08088_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08270_/B sky130_fd_sc_hd__xor2_1
XFILLER_107_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10050_ _15748_/Q _10057_/C _10009_/B vssd1 vssd1 vccd1 vccd1 _10050_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13740_ _13733_/C _13734_/C _13737_/Y _13738_/X vssd1 vssd1 vccd1 vccd1 _13741_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10952_ _15903_/Q _10992_/C _10951_/X vssd1 vssd1 vccd1 vccd1 _10954_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ _13696_/A _13671_/B _13671_/C vssd1 vssd1 vccd1 vccd1 _13672_/A sky130_fd_sc_hd__and3_1
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10883_ _10881_/A _10881_/B _10882_/X vssd1 vssd1 vccd1 vccd1 _15892_/D sky130_fd_sc_hd__a21oi_1
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15410_ _16157_/Q _16156_/Q _16155_/Q _15409_/X vssd1 vssd1 vccd1 vccd1 _16590_/D
+ sky130_fd_sc_hd__o31a_2
X_12622_ _16138_/Q _12622_/B _12628_/C vssd1 vssd1 vccd1 vccd1 _12622_/Y sky130_fd_sc_hd__nand3_1
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16390_ input11/X _16390_/D vssd1 vssd1 vccd1 vccd1 _16390_/Q sky130_fd_sc_hd__dfxtp_2
X_15341_ _16550_/Q _15341_/B _15346_/C vssd1 vssd1 vccd1 vccd1 _15348_/A sky130_fd_sc_hd__and3_1
X_12553_ _16130_/Q _12776_/B _12554_/C vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__and3_1
XFILLER_8_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11504_ _11617_/A _11509_/C vssd1 vssd1 vccd1 vccd1 _11504_/X sky130_fd_sc_hd__or2_1
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15272_ _15270_/A _15270_/B _15271_/X vssd1 vssd1 vccd1 vccd1 _16530_/D sky130_fd_sc_hd__a21oi_1
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ _12505_/A _12484_/B _12484_/C vssd1 vssd1 vccd1 vccd1 _12485_/A sky130_fd_sc_hd__and3_1
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14223_ _14237_/C vssd1 vssd1 vccd1 vccd1 _14245_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11435_ _15972_/Q _11444_/C _11434_/X vssd1 vssd1 vccd1 vccd1 _11435_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366_ _15963_/Q _11375_/C _11202_/X vssd1 vssd1 vccd1 vccd1 _11366_/Y sky130_fd_sc_hd__a21oi_1
X_14154_ _16357_/Q _14207_/B _14154_/C vssd1 vssd1 vccd1 vccd1 _14162_/B sky130_fd_sc_hd__and3_1
XFILLER_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10317_ _11384_/A vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13105_ _16208_/Q _13164_/B _13112_/C vssd1 vssd1 vccd1 vccd1 _13107_/C sky130_fd_sc_hd__nand3_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11297_ _11297_/A _11297_/B _11297_/C vssd1 vssd1 vccd1 vccd1 _11298_/C sky130_fd_sc_hd__nand3_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14085_ _16347_/Q _14193_/B _14094_/C vssd1 vssd1 vccd1 vccd1 _14085_/X sky130_fd_sc_hd__and3_1
XFILLER_125_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _10244_/Y _10247_/X _10240_/C _10241_/C vssd1 vssd1 vccd1 vccd1 _10250_/B
+ sky130_fd_sc_hd__o211ai_1
X_13036_ _13151_/A _13036_/B _13036_/C vssd1 vssd1 vccd1 vccd1 _13037_/C sky130_fd_sc_hd__or3_1
XFILLER_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10179_ _10179_/A _10179_/B _10186_/A vssd1 vssd1 vccd1 vccd1 _15769_/D sky130_fd_sc_hd__nor3_1
XFILLER_93_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14987_ _16484_/Q _14995_/C _14872_/X vssd1 vssd1 vccd1 vccd1 _14987_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16726_ _16726_/A _07830_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
XFILLER_47_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13938_ _13939_/B _13939_/C _13829_/X vssd1 vssd1 vccd1 vccd1 _13940_/B sky130_fd_sc_hd__o21ai_1
XFILLER_35_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13869_ _16316_/Q _13869_/B _13869_/C vssd1 vssd1 vccd1 vccd1 _13877_/A sky130_fd_sc_hd__and3_1
XFILLER_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15608_ _15812_/CLK _15608_/D vssd1 vssd1 vccd1 vccd1 _15608_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16588_ _16607_/CLK _16588_/D vssd1 vssd1 vccd1 vccd1 _16588_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_148_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _16551_/CLK _15539_/D vssd1 vssd1 vccd1 vccd1 _15539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ _09142_/A _09060_/B _09060_/C vssd1 vssd1 vccd1 vccd1 _09061_/A sky130_fd_sc_hd__and3_1
XFILLER_129_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ _16557_/Q _15885_/Q vssd1 vssd1 vccd1 vccd1 _08012_/C sky130_fd_sc_hd__or2_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09962_ _09962_/A _09962_/B vssd1 vssd1 vccd1 vccd1 _09962_/X sky130_fd_sc_hd__or2_1
X_08913_ _08911_/A _08911_/B _08912_/X vssd1 vssd1 vccd1 vccd1 _15511_/D sky130_fd_sc_hd__a21oi_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _15058_/A vssd1 vssd1 vccd1 vccd1 _10716_/A sky130_fd_sc_hd__clkbuf_2
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08844_ _15503_/Q _08866_/C _08843_/X vssd1 vssd1 vccd1 vccd1 _08846_/B sky130_fd_sc_hd__a21oi_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08775_ _08768_/C _08769_/C _08771_/Y _08781_/A vssd1 vssd1 vccd1 vccd1 _08781_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_27_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09327_ _09327_/A vssd1 vssd1 vccd1 vccd1 _15599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09258_ _15593_/Q _09267_/C _09992_/B vssd1 vssd1 vccd1 vccd1 _09261_/B sky130_fd_sc_hd__a21o_1
X_08209_ _14113_/A _07999_/B _08208_/X vssd1 vssd1 vccd1 vccd1 _08211_/B sky130_fd_sc_hd__o21a_1
X_09189_ _10789_/B vssd1 vssd1 vccd1 vccd1 _10922_/B sky130_fd_sc_hd__buf_2
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11220_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11226_/C sky130_fd_sc_hd__nor2_1
XFILLER_107_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11151_ _15932_/Q _11161_/C _11150_/X vssd1 vssd1 vccd1 vccd1 _11151_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10102_ _10100_/Y _10096_/C _10098_/Y _10108_/A vssd1 vssd1 vccd1 vccd1 _10108_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_122_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11082_ _11082_/A vssd1 vssd1 vccd1 vccd1 _15921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10033_ _10034_/B _10034_/C _10034_/A vssd1 vssd1 vccd1 vccd1 _10035_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14910_ _16472_/Q _14918_/C _14851_/X vssd1 vssd1 vccd1 vccd1 _14914_/B sky130_fd_sc_hd__a21o_1
XFILLER_102_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15890_ _16553_/Q _15890_/D vssd1 vssd1 vccd1 vccd1 _15890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14841_ _14841_/A vssd1 vssd1 vccd1 vccd1 _16459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16625__30 vssd1 vssd1 vccd1 vccd1 _16625__30/HI _16691_/A sky130_fd_sc_hd__conb_1
XFILLER_84_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14772_ _14772_/A _14772_/B vssd1 vssd1 vccd1 vccd1 _14774_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ _16050_/Q _11987_/C _11875_/X vssd1 vssd1 vccd1 vccd1 _11984_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16511_ _16607_/CLK _16511_/D vssd1 vssd1 vccd1 vccd1 _16511_/Q sky130_fd_sc_hd__dfxtp_1
X_13723_ _13759_/C vssd1 vssd1 vccd1 vccd1 _13765_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10935_ _10935_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__or2_1
XFILLER_140_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16442_ _16607_/CLK _16442_/D vssd1 vssd1 vccd1 vccd1 _16442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13654_ _13881_/A vssd1 vssd1 vccd1 vccd1 _13696_/A sky130_fd_sc_hd__clkbuf_2
X_10866_ _11150_/A vssd1 vssd1 vccd1 vccd1 _10866_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _12605_/A vssd1 vssd1 vccd1 vccd1 _12605_/X sky130_fd_sc_hd__clkbuf_4
X_16373_ _16389_/CLK _16373_/D vssd1 vssd1 vccd1 vccd1 _16373_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13585_ _16276_/Q _13592_/C _13414_/X vssd1 vssd1 vccd1 vccd1 _13585_/Y sky130_fd_sc_hd__a21oi_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ _15882_/Q _10797_/B _10805_/C vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__and3_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _15324_/A vssd1 vssd1 vccd1 vccd1 _15324_/Y sky130_fd_sc_hd__inv_2
X_12536_ _12653_/A _12536_/B _12540_/A vssd1 vssd1 vccd1 vccd1 _16126_/D sky130_fd_sc_hd__nor3_1
XFILLER_129_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15255_ _16528_/Q _15255_/B _15261_/C vssd1 vssd1 vccd1 vccd1 _15255_/Y sky130_fd_sc_hd__nand3_1
XFILLER_144_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ _12465_/A _12465_/B _12466_/X vssd1 vssd1 vccd1 vccd1 _16116_/D sky130_fd_sc_hd__a21oi_1
XFILLER_126_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14206_ _16365_/Q _14207_/C _13986_/X vssd1 vssd1 vccd1 vccd1 _14208_/A sky130_fd_sc_hd__a21oi_1
X_11418_ _12269_/A vssd1 vssd1 vccd1 vccd1 _11644_/B sky130_fd_sc_hd__clkbuf_2
X_15186_ _15186_/A vssd1 vssd1 vccd1 vccd1 _16516_/D sky130_fd_sc_hd__clkbuf_1
X_12398_ _12398_/A _12398_/B _12398_/C vssd1 vssd1 vccd1 vccd1 _12399_/A sky130_fd_sc_hd__and3_1
XFILLER_125_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14137_ _14135_/Y _14130_/C _14133_/Y _14134_/X vssd1 vssd1 vccd1 vccd1 _14138_/C
+ sky130_fd_sc_hd__a211o_1
X_11349_ _11349_/A _11349_/B _11349_/C vssd1 vssd1 vccd1 vccd1 _11350_/C sky130_fd_sc_hd__nand3_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14068_ _14068_/A _14068_/B _14068_/C vssd1 vssd1 vccd1 vccd1 _14069_/C sky130_fd_sc_hd__nand3_1
XFILLER_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13019_ _13019_/A _13019_/B _13019_/C vssd1 vssd1 vccd1 vccd1 _13020_/A sky130_fd_sc_hd__and3_1
XFILLER_66_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08560_ _08567_/A _08567_/B vssd1 vssd1 vccd1 vccd1 _15327_/A sky130_fd_sc_hd__xnor2_2
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08491_ _08477_/B _08491_/B vssd1 vssd1 vccd1 vccd1 _08532_/A sky130_fd_sc_hd__and2b_1
X_16709_ _16709_/A _07810_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_23_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09112_ _09112_/A _09112_/B vssd1 vssd1 vccd1 vccd1 _09114_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09043_ _08923_/X _09041_/A _09039_/X vssd1 vssd1 vccd1 vccd1 _09044_/B sky130_fd_sc_hd__o21ai_1
XFILLER_136_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09945_ _15727_/Q _09945_/B _09945_/C vssd1 vssd1 vccd1 vccd1 _09950_/A sky130_fd_sc_hd__and3_1
XFILLER_131_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09946_/A _09876_/B _09879_/B vssd1 vssd1 vccd1 vccd1 _15708_/D sky130_fd_sc_hd__nor3_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08825_/A _08825_/B _08826_/X vssd1 vssd1 vccd1 vccd1 _15493_/D sky130_fd_sc_hd__a21oi_1
XFILLER_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _08854_/A vssd1 vssd1 vccd1 vccd1 _08846_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _15470_/Q _09271_/A _08689_/C vssd1 vssd1 vccd1 vccd1 _08690_/B sky130_fd_sc_hd__and3_1
XFILLER_14_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _15857_/Q _15856_/Q _15855_/Q _10719_/X vssd1 vssd1 vccd1 vccd1 _15867_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10651_ _15856_/Q _10658_/C _10454_/X vssd1 vssd1 vccd1 vccd1 _10651_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10582_ _15843_/Q _10612_/C _10426_/X vssd1 vssd1 vccd1 vccd1 _10584_/B sky130_fd_sc_hd__a21oi_1
X_13370_ _13368_/A _13368_/B _13369_/X vssd1 vssd1 vccd1 vccd1 _16244_/D sky130_fd_sc_hd__a21oi_1
X_12321_ _12343_/A _12321_/B _12321_/C vssd1 vssd1 vccd1 vccd1 _12322_/A sky130_fd_sc_hd__and3_1
XFILLER_126_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15040_ _16493_/Q _15049_/C _14872_/X vssd1 vssd1 vccd1 vccd1 _15040_/Y sky130_fd_sc_hd__a21oi_1
X_12252_ _16087_/Q _12252_/B _12263_/C vssd1 vssd1 vccd1 vccd1 _12257_/A sky130_fd_sc_hd__and3_1
XFILLER_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11203_ _15939_/Q _11211_/C _11202_/X vssd1 vssd1 vccd1 vccd1 _11203_/Y sky130_fd_sc_hd__a21oi_1
X_12183_ _12183_/A _12187_/C vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__or2_1
XFILLER_122_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ input3/X vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__buf_2
XFILLER_96_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15942_ _15365_/A _15942_/D vssd1 vssd1 vccd1 vccd1 _15942_/Q sky130_fd_sc_hd__dfxtp_2
X_11065_ _11066_/B _11066_/C _11066_/A vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__a21o_1
XFILLER_1_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10016_ _10016_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _10017_/B sky130_fd_sc_hd__and2_1
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15873_ _16570_/CLK _15873_/D vssd1 vssd1 vccd1 vccd1 _15873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14824_ _16457_/Q _14882_/B _14831_/C vssd1 vssd1 vccd1 vccd1 _14824_/Y sky130_fd_sc_hd__nand3_1
XFILLER_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14755_ _16448_/Q _14764_/C _14588_/X vssd1 vssd1 vccd1 vccd1 _14755_/Y sky130_fd_sc_hd__a21oi_1
X_11967_ _12002_/C vssd1 vssd1 vccd1 vccd1 _12010_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13706_ _16293_/Q _13709_/C _13705_/X vssd1 vssd1 vccd1 vccd1 _13710_/A sky130_fd_sc_hd__a21oi_1
X_10918_ _10918_/A vssd1 vssd1 vccd1 vccd1 _15897_/D sky130_fd_sc_hd__clkbuf_1
X_14686_ _14707_/A _14686_/B _14686_/C vssd1 vssd1 vccd1 vccd1 _14687_/A sky130_fd_sc_hd__and3_1
XFILLER_60_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11898_ _11898_/A _11905_/B vssd1 vssd1 vccd1 vccd1 _11900_/A sky130_fd_sc_hd__or2_1
X_16425_ _16595_/CLK _16425_/D vssd1 vssd1 vccd1 vccd1 _16425_/Q sky130_fd_sc_hd__dfxtp_2
X_13637_ _16284_/Q _13645_/C _13414_/X vssd1 vssd1 vccd1 vccd1 _13637_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10849_ _15890_/Q _10852_/C _14932_/A vssd1 vssd1 vccd1 vccd1 _10849_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16356_ _16389_/CLK _16356_/D vssd1 vssd1 vccd1 vccd1 _16356_/Q sky130_fd_sc_hd__dfxtp_1
X_13568_ _13583_/A _13568_/B _13568_/C vssd1 vssd1 vccd1 vccd1 _13569_/A sky130_fd_sc_hd__and3_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ _16709_/A _15321_/B _15307_/C vssd1 vssd1 vccd1 vccd1 _15324_/A sky130_fd_sc_hd__and3_1
X_12519_ _12801_/A vssd1 vssd1 vccd1 vccd1 _12749_/A sky130_fd_sc_hd__clkbuf_2
X_16287_ _16533_/Q _16287_/D vssd1 vssd1 vccd1 vccd1 _16287_/Q sky130_fd_sc_hd__dfxtp_1
X_13499_ _16264_/Q _13507_/C _13443_/X vssd1 vssd1 vccd1 vccd1 _13503_/B sky130_fd_sc_hd__a21o_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15238_ _15258_/A _15238_/B _15238_/C vssd1 vssd1 vccd1 vccd1 _15239_/A sky130_fd_sc_hd__and3_1
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _15274_/A _15169_/B _15169_/C vssd1 vssd1 vccd1 vccd1 _15170_/C sky130_fd_sc_hd__or3_1
XFILLER_114_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07991_ _16571_/Q _07991_/B _08204_/A vssd1 vssd1 vccd1 vccd1 _08204_/B sky130_fd_sc_hd__nand3_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09730_ _09841_/A _09730_/B _09733_/B vssd1 vssd1 vccd1 vccd1 _15681_/D sky130_fd_sc_hd__nor3_1
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ _09615_/X _09656_/B _09572_/X vssd1 vssd1 vccd1 vccd1 _09663_/A sky130_fd_sc_hd__a21oi_1
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08612_ input3/X vssd1 vssd1 vccd1 vccd1 _13288_/A sky130_fd_sc_hd__buf_2
X_09592_ _15657_/Q _09636_/B _09592_/C vssd1 vssd1 vccd1 vccd1 _09598_/A sky130_fd_sc_hd__and3_1
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08543_ _08543_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _08556_/B sky130_fd_sc_hd__xor2_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08474_ _08407_/A _08407_/B _08473_/Y vssd1 vssd1 vccd1 vccd1 _08475_/B sky130_fd_sc_hd__a21oi_2
XFILLER_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09026_ _15542_/Q _09028_/C _08989_/X vssd1 vssd1 vccd1 vccd1 _09029_/A sky130_fd_sc_hd__a21oi_1
XFILLER_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09928_ _09924_/Y _09927_/X _09894_/X vssd1 vssd1 vccd1 vccd1 _09928_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_120_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09859_ _09953_/A vssd1 vssd1 vccd1 vccd1 _09946_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12870_ _12870_/A vssd1 vssd1 vccd1 vccd1 _16173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _16025_/Q _11878_/B _11821_/C vssd1 vssd1 vccd1 vccd1 _11821_/Y sky130_fd_sc_hd__nand3_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _16412_/Q _14598_/B _14547_/C vssd1 vssd1 vccd1 vccd1 _14540_/Y sky130_fd_sc_hd__nand3_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11752_/A _11752_/B _11752_/C vssd1 vssd1 vccd1 vccd1 _11753_/C sky130_fd_sc_hd__nand3_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10699_/Y _10709_/A _10702_/Y _10695_/C vssd1 vssd1 vccd1 vccd1 _10705_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _16403_/Q _14480_/C _14308_/X vssd1 vssd1 vccd1 vccd1 _14471_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11683_/A vssd1 vssd1 vccd1 vccd1 _11698_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16237_/CLK _16210_/D vssd1 vssd1 vccd1 vccd1 _16210_/Q sky130_fd_sc_hd__dfxtp_1
X_13422_ _16253_/Q _13424_/C _13421_/X vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__a21oi_1
X_10634_ _10635_/B _10635_/C _10635_/A vssd1 vssd1 vccd1 vccd1 _10636_/B sky130_fd_sc_hd__a21o_1
X_16141_ _16555_/Q _16141_/D vssd1 vssd1 vccd1 vccd1 _16141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353_ _13351_/Y _13347_/C _13349_/Y _13350_/X vssd1 vssd1 vccd1 vccd1 _13354_/C
+ sky130_fd_sc_hd__a211o_1
X_10565_ _15839_/Q _10707_/B _10565_/C vssd1 vssd1 vccd1 vccd1 _10566_/B sky130_fd_sc_hd__and3_1
XFILLER_127_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _12304_/A _12304_/B _12304_/C vssd1 vssd1 vccd1 vccd1 _12305_/C sky130_fd_sc_hd__or3_1
X_16072_ _16118_/CLK _16072_/D vssd1 vssd1 vccd1 vccd1 _16072_/Q sky130_fd_sc_hd__dfxtp_1
X_13284_ _13282_/Y _13283_/X _13279_/C _13280_/C vssd1 vssd1 vccd1 vccd1 _13286_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_6_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10496_ _10489_/C _10490_/C _10493_/Y _10494_/X vssd1 vssd1 vccd1 vccd1 _10497_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15023_ _15023_/A _15023_/B _15023_/C vssd1 vssd1 vccd1 vccd1 _15024_/C sky130_fd_sc_hd__nand3_1
X_12235_ _12801_/A vssd1 vssd1 vccd1 vccd1 _12466_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12166_ _16075_/Q _12218_/B _12173_/C vssd1 vssd1 vccd1 vccd1 _12166_/X sky130_fd_sc_hd__and3_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11117_ _15927_/Q _11161_/C _10951_/X vssd1 vssd1 vccd1 vccd1 _11119_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12097_ _12097_/A vssd1 vssd1 vccd1 vccd1 _16064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15925_ _15365_/A _15925_/D vssd1 vssd1 vccd1 vccd1 _15925_/Q sky130_fd_sc_hd__dfxtp_1
X_11048_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11053_/C sky130_fd_sc_hd__nor2_1
XFILLER_110_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 io_in[26] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_6
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ _16570_/CLK _15856_/D vssd1 vssd1 vccd1 vccd1 _15856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14807_ _16456_/Q _15033_/B _14808_/C vssd1 vssd1 vccd1 vccd1 _14807_/X sky130_fd_sc_hd__and3_1
X_15787_ _15791_/CLK _15787_/D vssd1 vssd1 vccd1 vccd1 _15787_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ _12999_/A vssd1 vssd1 vccd1 vccd1 _16191_/D sky130_fd_sc_hd__clkbuf_1
X_14738_ _14738_/A _14738_/B _14738_/C vssd1 vssd1 vccd1 vccd1 _14739_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14669_ _14669_/A vssd1 vssd1 vccd1 vccd1 _14669_/X sky130_fd_sc_hd__clkbuf_2
X_16408_ input11/X _16408_/D vssd1 vssd1 vccd1 vccd1 _16408_/Q sky130_fd_sc_hd__dfxtp_1
X_08190_ _08190_/A _08190_/B vssd1 vssd1 vccd1 vccd1 _08346_/A sky130_fd_sc_hd__xnor2_4
X_16339_ _16346_/CLK _16339_/D vssd1 vssd1 vccd1 vccd1 _16339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07974_ _09541_/C _07974_/B vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__xnor2_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09713_ _09727_/C vssd1 vssd1 vccd1 vccd1 _09739_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09644_ _10112_/A vssd1 vssd1 vccd1 vccd1 _09644_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09575_ _09575_/A _09575_/B vssd1 vssd1 vccd1 vccd1 _15650_/D sky130_fd_sc_hd__nor2_1
XFILLER_70_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _08526_/A vssd1 vssd1 vccd1 vccd1 _10430_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08457_ _08497_/A _08497_/B vssd1 vssd1 vccd1 vccd1 _08462_/A sky130_fd_sc_hd__xor2_1
X_08388_ _08388_/A _08388_/B vssd1 vssd1 vccd1 vccd1 _08388_/X sky130_fd_sc_hd__or2_1
XFILLER_136_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _10347_/Y _10348_/X _10349_/Y _10345_/C vssd1 vssd1 vccd1 vccd1 _10352_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_137_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09009_ _15524_/Q _15523_/Q _15522_/Q _08887_/X vssd1 vssd1 vccd1 vccd1 _15534_/D
+ sky130_fd_sc_hd__o31a_1
X_10281_ _10285_/B vssd1 vssd1 vccd1 vccd1 _10294_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ _12020_/A vssd1 vssd1 vccd1 vccd1 _16053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13971_ _16331_/Q _13981_/C _13750_/X vssd1 vssd1 vccd1 vccd1 _13971_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15710_ _15812_/CLK _15710_/D vssd1 vssd1 vccd1 vccd1 _15710_/Q sky130_fd_sc_hd__dfxtp_1
X_12922_ _13034_/A vssd1 vssd1 vccd1 vccd1 _12963_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16690_ _16690_/A _07787_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ _15812_/CLK _15641_/D vssd1 vssd1 vccd1 vccd1 _15641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ _16171_/Q _12911_/B _12860_/C vssd1 vssd1 vccd1 vccd1 _12853_/Y sky130_fd_sc_hd__nand3_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _16023_/Q _11969_/B _11814_/C vssd1 vssd1 vccd1 vccd1 _11810_/A sky130_fd_sc_hd__and3_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15812_/CLK _15572_/D vssd1 vssd1 vccd1 vccd1 _15572_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _16163_/Q _12784_/B _12792_/C vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__and3_1
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _16411_/Q _14748_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _14523_/X sky130_fd_sc_hd__and3_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11735_ _11903_/A vssd1 vssd1 vccd1 vccd1 _11776_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14454_ _14454_/A _14454_/B _14454_/C vssd1 vssd1 vccd1 vccd1 _14455_/C sky130_fd_sc_hd__nand3_1
X_11666_ _11666_/A _11666_/B _11670_/B vssd1 vssd1 vccd1 vccd1 _16003_/D sky130_fd_sc_hd__nor3_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13405_ _13405_/A vssd1 vssd1 vccd1 vccd1 _16249_/D sky130_fd_sc_hd__clkbuf_1
X_10617_ _10615_/A _10615_/B _10616_/X vssd1 vssd1 vccd1 vccd1 _15846_/D sky130_fd_sc_hd__a21oi_1
X_14385_ _14383_/A _14383_/B _14384_/X vssd1 vssd1 vccd1 vccd1 _16388_/D sky130_fd_sc_hd__a21oi_1
X_11597_ _11604_/A _11597_/B _11597_/C vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__and3_1
XFILLER_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ _16554_/Q _16124_/D vssd1 vssd1 vccd1 vccd1 _16124_/Q sky130_fd_sc_hd__dfxtp_1
X_13336_ _16241_/Q _13336_/B _13336_/C vssd1 vssd1 vccd1 vccd1 _13336_/X sky130_fd_sc_hd__and3_1
X_10548_ _10541_/C _10542_/C _10544_/Y _10546_/X vssd1 vssd1 vccd1 vccd1 _10549_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ _16118_/CLK _16055_/D vssd1 vssd1 vccd1 vccd1 _16055_/Q sky130_fd_sc_hd__dfxtp_1
X_13267_ _13302_/A _13267_/B _13267_/C vssd1 vssd1 vccd1 vccd1 _13268_/A sky130_fd_sc_hd__and3_1
X_10479_ _10483_/C vssd1 vssd1 vccd1 vccd1 _10494_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15006_ _15004_/A _15004_/B _15005_/X vssd1 vssd1 vccd1 vccd1 _16485_/D sky130_fd_sc_hd__a21oi_1
X_12218_ _16083_/Q _12218_/B _12226_/C vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__and3_1
X_13198_ _16221_/Q _13199_/C _13140_/X vssd1 vssd1 vccd1 vccd1 _13200_/A sky130_fd_sc_hd__a21oi_1
XFILLER_2_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12149_ _12170_/A _12149_/B _12149_/C vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__and3_1
XFILLER_123_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15908_ _16553_/Q _15908_/D vssd1 vssd1 vccd1 vccd1 _15908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15839_ _16551_/CLK _15839_/D vssd1 vssd1 vccd1 vccd1 _15839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09360_ _15610_/Q _09448_/B _09360_/C vssd1 vssd1 vccd1 vccd1 _09366_/A sky130_fd_sc_hd__and3_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08311_ _15350_/A vssd1 vssd1 vccd1 vccd1 _15344_/A sky130_fd_sc_hd__buf_2
X_09291_ _09744_/A vssd1 vssd1 vccd1 vccd1 _09291_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _08380_/A _08380_/B vssd1 vssd1 vccd1 vccd1 _08370_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_24 _10016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _13392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ _07933_/A _07933_/B _07945_/B _07944_/B _11798_/A vssd1 vssd1 vccd1 vccd1
+ _08328_/B sky130_fd_sc_hd__o32a_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07957_ _07957_/A _07957_/B vssd1 vssd1 vccd1 vccd1 _07958_/B sky130_fd_sc_hd__nand2_2
XFILLER_56_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07888_ _14279_/A _07888_/B vssd1 vssd1 vccd1 vccd1 _07889_/B sky130_fd_sc_hd__xnor2_4
XFILLER_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _09812_/A vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09558_ _09557_/X _09556_/Y _09424_/X vssd1 vssd1 vccd1 vccd1 _09558_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08509_ _08509_/A _08509_/B _08509_/C vssd1 vssd1 vccd1 vccd1 _08510_/B sky130_fd_sc_hd__and3_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09489_ _09489_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _15632_/D sky130_fd_sc_hd__nor2_1
XFILLER_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11520_ _11520_/A _11520_/B _11525_/A vssd1 vssd1 vccd1 vccd1 _15982_/D sky130_fd_sc_hd__nor3_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ _11452_/B _11452_/C _11282_/X vssd1 vssd1 vccd1 vccd1 _11453_/B sky130_fd_sc_hd__o21ai_1
X_10402_ _15811_/Q _10402_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10410_/A sky130_fd_sc_hd__and3_1
X_14170_ _16359_/Q _14227_/B _14179_/C vssd1 vssd1 vccd1 vccd1 _14175_/A sky130_fd_sc_hd__and3_1
X_11382_ _11382_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__or2_1
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ _13117_/Y _13119_/X _13120_/Y _13115_/C vssd1 vssd1 vccd1 vccd1 _13123_/B
+ sky130_fd_sc_hd__o211ai_1
X_10333_ _10429_/A _10333_/B _10337_/A vssd1 vssd1 vccd1 vccd1 _15796_/D sky130_fd_sc_hd__nor3_1
X_13052_ _16201_/Q _13062_/C _12887_/X vssd1 vssd1 vccd1 vccd1 _13052_/Y sky130_fd_sc_hd__a21oi_1
X_10264_ _10262_/Y _10258_/C _10260_/Y _10269_/A vssd1 vssd1 vccd1 vccd1 _10269_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_87_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12003_ _16051_/Q _12060_/B _12010_/C vssd1 vssd1 vccd1 vccd1 _12003_/Y sky130_fd_sc_hd__nand3_1
X_10195_ _15774_/Q _10206_/C _10138_/X vssd1 vssd1 vccd1 vccd1 _10195_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16742_ _16742_/A _07758_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
X_13954_ _13977_/A _13954_/B _13954_/C vssd1 vssd1 vccd1 vccd1 _13955_/A sky130_fd_sc_hd__and3_1
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12905_ _12902_/Y _12903_/X _12904_/Y _12899_/C vssd1 vssd1 vccd1 vccd1 _12907_/B
+ sky130_fd_sc_hd__o211ai_1
X_13885_ _13885_/A vssd1 vssd1 vccd1 vccd1 _16317_/D sky130_fd_sc_hd__clkbuf_1
X_16670__75 vssd1 vssd1 vccd1 vccd1 _16670__75/HI _16746_/A sky130_fd_sc_hd__conb_1
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15624_ _16551_/CLK _15624_/D vssd1 vssd1 vccd1 vccd1 _15624_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ _16169_/Q _13009_/B _12836_/C vssd1 vssd1 vccd1 vccd1 _12836_/Y sky130_fd_sc_hd__nand3_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15555_ _15791_/CLK _15555_/D vssd1 vssd1 vccd1 vccd1 _15555_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12788_/A _12767_/B _12767_/C vssd1 vssd1 vccd1 vccd1 _12768_/A sky130_fd_sc_hd__and3_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _16408_/Q _14506_/B _14516_/C vssd1 vssd1 vccd1 vccd1 _14511_/A sky130_fd_sc_hd__and3_1
XFILLER_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11718_ _11718_/A vssd1 vssd1 vccd1 vccd1 _16010_/D sky130_fd_sc_hd__clkbuf_1
X_15486_ _16570_/CLK _15486_/D vssd1 vssd1 vccd1 vccd1 _15486_/Q sky130_fd_sc_hd__dfxtp_1
X_12698_ _12751_/A vssd1 vssd1 vccd1 vccd1 _12736_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14437_ _14437_/A _14441_/C vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__or2_1
X_11649_ _11643_/Y _11644_/X _11648_/Y _11641_/C vssd1 vssd1 vccd1 vccd1 _11651_/B
+ sky130_fd_sc_hd__o211ai_1
Xinput11 wb_clk_i vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_12
X_14368_ _14366_/Y _14361_/C _14363_/Y _14364_/X vssd1 vssd1 vccd1 vccd1 _14369_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16107_ _16118_/CLK _16107_/D vssd1 vssd1 vccd1 vccd1 _16107_/Q sky130_fd_sc_hd__dfxtp_1
X_13319_ _13432_/A _13319_/B _13319_/C vssd1 vssd1 vccd1 vccd1 _13320_/C sky130_fd_sc_hd__or3_1
XFILLER_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14299_ _14314_/A _14299_/B _14299_/C vssd1 vssd1 vccd1 vccd1 _14300_/A sky130_fd_sc_hd__and3_1
XFILLER_143_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16038_ _16118_/CLK _16038_/D vssd1 vssd1 vccd1 vccd1 _16038_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08860_ _15505_/Q _08866_/C _08859_/X vssd1 vssd1 vccd1 vccd1 _08860_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07811_ _07811_/A vssd1 vssd1 vccd1 vccd1 _07811_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08791_ _08921_/A _08921_/B _08791_/C vssd1 vssd1 vccd1 vccd1 _08793_/A sky130_fd_sc_hd__and3_1
XFILLER_38_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09412_ _09412_/A _09412_/B _09412_/C vssd1 vssd1 vccd1 vccd1 _09413_/C sky130_fd_sc_hd__nand3_1
XFILLER_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09343_ _09339_/Y _09342_/X _09304_/X vssd1 vssd1 vccd1 vccd1 _09343_/Y sky130_fd_sc_hd__a21oi_1
X_09274_ _15255_/B vssd1 vssd1 vccd1 vccd1 _09837_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08225_ _08225_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08226_/B sky130_fd_sc_hd__xor2_2
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08156_ _08157_/A _08157_/B vssd1 vssd1 vccd1 vccd1 _08353_/A sky130_fd_sc_hd__nand2_2
XFILLER_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08087_ _15121_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08088_/B sky130_fd_sc_hd__xnor2_2
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08989_ _15346_/B vssd1 vssd1 vccd1 vccd1 _08989_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10951_ _11233_/A vssd1 vssd1 vccd1 vccd1 _10951_/X sky130_fd_sc_hd__buf_2
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13670_ _13670_/A _13670_/B _13670_/C vssd1 vssd1 vccd1 vccd1 _13671_/C sky130_fd_sc_hd__nand3_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10882_ _11049_/A _10886_/C vssd1 vssd1 vccd1 vccd1 _10882_/X sky130_fd_sc_hd__or2_1
XFILLER_71_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12621_ _16139_/Q _12784_/B _12628_/C vssd1 vssd1 vccd1 vccd1 _12621_/X sky130_fd_sc_hd__and3_1
X_15340_ _16550_/Q _15346_/C _10301_/C vssd1 vssd1 vccd1 vccd1 _15340_/Y sky130_fd_sc_hd__a21oi_1
X_12552_ _13682_/A vssd1 vssd1 vccd1 vccd1 _12776_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ _11503_/A _11503_/B vssd1 vssd1 vccd1 vccd1 _11509_/C sky130_fd_sc_hd__nor2_1
X_15271_ _15271_/A _15274_/C vssd1 vssd1 vccd1 vccd1 _15271_/X sky130_fd_sc_hd__or2_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12483_ _12483_/A _12483_/B _12483_/C vssd1 vssd1 vccd1 vccd1 _12484_/C sky130_fd_sc_hd__nand3_1
XFILLER_138_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14222_ _14222_/A vssd1 vssd1 vccd1 vccd1 _14237_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11434_ _12567_/A vssd1 vssd1 vccd1 vccd1 _11434_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14153_ _16357_/Q _14154_/C _13986_/X vssd1 vssd1 vccd1 vccd1 _14155_/A sky130_fd_sc_hd__a21oi_1
X_11365_ _11365_/A vssd1 vssd1 vccd1 vccd1 _15961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13104_ _16208_/Q _13112_/C _12879_/X vssd1 vssd1 vccd1 vccd1 _13107_/B sky130_fd_sc_hd__a21o_1
XFILLER_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10316_ _13085_/A vssd1 vssd1 vccd1 vccd1 _11384_/A sky130_fd_sc_hd__buf_4
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14084_ _16347_/Q _14094_/C _14029_/X vssd1 vssd1 vccd1 vccd1 _14084_/Y sky130_fd_sc_hd__a21oi_1
X_11296_ _11297_/B _11297_/C _11297_/A vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__a21o_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _13036_/B _13036_/C _12982_/X vssd1 vssd1 vccd1 vccd1 _13037_/B sky130_fd_sc_hd__o21ai_1
XFILLER_140_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10247_ _15782_/Q _10494_/B _10247_/C vssd1 vssd1 vccd1 vccd1 _10247_/X sky130_fd_sc_hd__and3_1
XFILLER_79_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10178_ _15771_/Q _10178_/B _10178_/C vssd1 vssd1 vccd1 vccd1 _10186_/A sky130_fd_sc_hd__and3_1
XFILLER_94_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14986_ _14986_/A vssd1 vssd1 vccd1 vccd1 _16482_/D sky130_fd_sc_hd__clkbuf_1
X_16725_ _16725_/A _07829_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13937_ _14160_/A vssd1 vssd1 vccd1 vccd1 _13977_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13868_ _16316_/Q _13875_/C _13698_/X vssd1 vssd1 vccd1 vccd1 _13868_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15607_ _16551_/CLK _15607_/D vssd1 vssd1 vccd1 vccd1 _15607_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ _12936_/A _12819_/B _12823_/A vssd1 vssd1 vccd1 vccd1 _16166_/D sky130_fd_sc_hd__nor3_1
XFILLER_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16587_ _16607_/CLK _16587_/D vssd1 vssd1 vccd1 vccd1 _16587_/Q sky130_fd_sc_hd__dfxtp_1
X_13799_ _16306_/Q _13906_/B _13800_/C vssd1 vssd1 vccd1 vccd1 _13799_/X sky130_fd_sc_hd__and3_1
X_15538_ _16551_/CLK _15538_/D vssd1 vssd1 vccd1 vccd1 _15538_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15469_ _16551_/CLK _15469_/D vssd1 vssd1 vccd1 vccd1 _15469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08010_ _16557_/Q _15885_/Q vssd1 vssd1 vccd1 vccd1 _08218_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09961_ _09961_/A _09961_/B vssd1 vssd1 vccd1 vccd1 _09961_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08912_ _09074_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _08912_/X sky130_fd_sc_hd__or2_1
X_09892_ _09744_/X _09890_/B _09891_/Y vssd1 vssd1 vccd1 vccd1 _15711_/D sky130_fd_sc_hd__o21a_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _08843_/A vssd1 vssd1 vccd1 vccd1 _08843_/X sky130_fd_sc_hd__clkbuf_4
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08774_ _08771_/Y _08781_/A _08768_/C _08769_/C vssd1 vssd1 vccd1 vccd1 _08776_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09326_ _09367_/A _09326_/B _09326_/C vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__and3_1
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ _10183_/A vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__buf_2
X_08208_ _08208_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _08208_/X sky130_fd_sc_hd__or2_1
X_09188_ _09256_/A _09188_/B _09194_/B vssd1 vssd1 vccd1 vccd1 _15573_/D sky130_fd_sc_hd__nor3_1
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08139_ _08139_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08321_/A sky130_fd_sc_hd__xnor2_1
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ _11150_/A vssd1 vssd1 vccd1 vccd1 _11150_/X sky130_fd_sc_hd__buf_2
X_10101_ _10098_/Y _10108_/A _10100_/Y _10096_/C vssd1 vssd1 vccd1 vccd1 _10103_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11081_ _11088_/A _11081_/B _11081_/C vssd1 vssd1 vccd1 vccd1 _11082_/A sky130_fd_sc_hd__and3_1
XFILLER_68_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10032_ _15745_/Q _10288_/C _10038_/C vssd1 vssd1 vccd1 vccd1 _10034_/C sky130_fd_sc_hd__nand3_1
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14840_ _14878_/A _14840_/B _14840_/C vssd1 vssd1 vccd1 vccd1 _14841_/A sky130_fd_sc_hd__and3_1
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14771_ _14771_/A _14780_/B vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__or2_1
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11983_ _11983_/A vssd1 vssd1 vccd1 vccd1 _16048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16510_ _16607_/CLK _16510_/D vssd1 vssd1 vccd1 vccd1 _16510_/Q sky130_fd_sc_hd__dfxtp_1
X_13722_ _13745_/C vssd1 vssd1 vccd1 vccd1 _13759_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10934_ _15901_/Q _11099_/B _10934_/C vssd1 vssd1 vccd1 vccd1 _10944_/B sky130_fd_sc_hd__and3_1
X_16640__45 vssd1 vssd1 vccd1 vccd1 _16640__45/HI _16716_/A sky130_fd_sc_hd__conb_1
X_16441_ _16595_/CLK _16441_/D vssd1 vssd1 vccd1 vccd1 _16441_/Q sky130_fd_sc_hd__dfxtp_1
X_13653_ _14777_/A vssd1 vssd1 vccd1 vccd1 _13881_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10865_ _10865_/A vssd1 vssd1 vccd1 vccd1 _15890_/D sky130_fd_sc_hd__clkbuf_1
X_12604_ _12604_/A vssd1 vssd1 vccd1 vccd1 _16135_/D sky130_fd_sc_hd__clkbuf_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _16389_/CLK _16372_/D vssd1 vssd1 vccd1 vccd1 _16372_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _13584_/A vssd1 vssd1 vccd1 vccd1 _16274_/D sky130_fd_sc_hd__clkbuf_1
X_10796_ _15882_/Q _10805_/C _10456_/A vssd1 vssd1 vccd1 vccd1 _10796_/Y sky130_fd_sc_hd__a21oi_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15323_ _15320_/Y _15317_/Y _15322_/Y _15316_/B vssd1 vssd1 vccd1 vccd1 _15326_/B
+ sky130_fd_sc_hd__o211a_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _16127_/Q _12535_/B _12545_/C vssd1 vssd1 vccd1 vccd1 _12540_/A sky130_fd_sc_hd__and3_1
XFILLER_8_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15254_ _16529_/Q _15254_/B _15261_/C vssd1 vssd1 vccd1 vccd1 _15254_/X sky130_fd_sc_hd__and3_1
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12466_ _12466_/A _12470_/C vssd1 vssd1 vccd1 vccd1 _12466_/X sky130_fd_sc_hd__or2_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14205_ _14205_/A _14205_/B _14209_/B vssd1 vssd1 vccd1 vccd1 _16363_/D sky130_fd_sc_hd__nor3_1
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ _15970_/Q _11420_/C _11306_/X vssd1 vssd1 vccd1 vccd1 _11417_/Y sky130_fd_sc_hd__a21oi_1
X_15185_ _15205_/A _15185_/B _15185_/C vssd1 vssd1 vccd1 vccd1 _15186_/A sky130_fd_sc_hd__and3_1
X_12397_ _12395_/Y _12390_/C _12392_/Y _12393_/X vssd1 vssd1 vccd1 vccd1 _12398_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14136_ _14133_/Y _14134_/X _14135_/Y _14130_/C vssd1 vssd1 vccd1 vccd1 _14138_/B
+ sky130_fd_sc_hd__o211ai_1
X_11348_ _11349_/B _11349_/C _11349_/A vssd1 vssd1 vccd1 vccd1 _11350_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ _14068_/B _14068_/C _14068_/A vssd1 vssd1 vccd1 vccd1 _14069_/B sky130_fd_sc_hd__a21o_1
X_11279_ _11332_/A _11284_/C vssd1 vssd1 vccd1 vccd1 _11279_/X sky130_fd_sc_hd__or2_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13018_ _13016_/Y _13012_/C _13014_/Y _13015_/X vssd1 vssd1 vccd1 vccd1 _13019_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14969_ _14970_/B _14970_/C _14970_/A vssd1 vssd1 vccd1 vccd1 _14971_/B sky130_fd_sc_hd__a21o_1
X_16708_ _16708_/A _07809_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
X_08490_ _08490_/A vssd1 vssd1 vccd1 vccd1 _08561_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09111_ _09111_/A _09111_/B vssd1 vssd1 vccd1 vccd1 _09114_/A sky130_fd_sc_hd__or2_1
XFILLER_148_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09042_ _09124_/A _09124_/B _09042_/C vssd1 vssd1 vccd1 vccd1 _09044_/A sky130_fd_sc_hd__and3_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09944_ _15727_/Q _09966_/C _09943_/X vssd1 vssd1 vccd1 vccd1 _09946_/B sky130_fd_sc_hd__a21oi_1
XFILLER_131_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09875_ _09869_/C _09870_/C _09872_/Y _09879_/A vssd1 vssd1 vccd1 vccd1 _09879_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08870_/A _08826_/B vssd1 vssd1 vccd1 vccd1 _08826_/X sky130_fd_sc_hd__or2_1
XFILLER_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08757_ _15470_/Q _15469_/Q _15468_/Q _08667_/X vssd1 vssd1 vccd1 vccd1 _15480_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_39_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _15470_/Q _08689_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _08690_/A sky130_fd_sc_hd__a21oi_1
XFILLER_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10650_ _10650_/A vssd1 vssd1 vccd1 vccd1 _15853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ _09307_/X _09296_/B _09308_/X vssd1 vssd1 vccd1 vccd1 _09313_/A sky130_fd_sc_hd__a21oi_1
XFILLER_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10581_ _10606_/C vssd1 vssd1 vccd1 vccd1 _10612_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _12320_/A _12320_/B _12320_/C vssd1 vssd1 vccd1 vccd1 _12321_/C sky130_fd_sc_hd__nand3_1
X_12251_ _16087_/Q _12296_/C _12081_/X vssd1 vssd1 vccd1 vccd1 _12253_/B sky130_fd_sc_hd__a21oi_1
XFILLER_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ _12968_/A vssd1 vssd1 vccd1 vccd1 _11202_/X sky130_fd_sc_hd__buf_2
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _12182_/A _12182_/B vssd1 vssd1 vccd1 vccd1 _12187_/C sky130_fd_sc_hd__nor2_1
XFILLER_134_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11133_ _15930_/Q _11137_/C _11023_/X vssd1 vssd1 vccd1 vccd1 _11133_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15941_ _15365_/A _15941_/D vssd1 vssd1 vccd1 vccd1 _15941_/Q sky130_fd_sc_hd__dfxtp_1
X_11064_ _15920_/Q _11183_/B _11070_/C vssd1 vssd1 vccd1 vccd1 _11066_/C sky130_fd_sc_hd__nand3_1
XFILLER_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10015_ _10008_/Y _10009_/X _10011_/B vssd1 vssd1 vccd1 vccd1 _10016_/B sky130_fd_sc_hd__o21a_1
X_15872_ _16570_/CLK _15872_/D vssd1 vssd1 vccd1 vccd1 _15872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14823_ _16458_/Q _14995_/B _14823_/C vssd1 vssd1 vccd1 vccd1 _14833_/A sky130_fd_sc_hd__and3_1
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11966_ _11987_/C vssd1 vssd1 vccd1 vccd1 _12002_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14754_ _14754_/A vssd1 vssd1 vccd1 vccd1 _16446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _10925_/A _10917_/B _10917_/C vssd1 vssd1 vccd1 vccd1 _10918_/A sky130_fd_sc_hd__and3_1
X_13705_ _13705_/A vssd1 vssd1 vccd1 vccd1 _13705_/X sky130_fd_sc_hd__clkbuf_2
X_14685_ _14685_/A _14685_/B _14685_/C vssd1 vssd1 vccd1 vccd1 _14686_/C sky130_fd_sc_hd__nand3_1
X_11897_ _16037_/Q _11950_/B _11897_/C vssd1 vssd1 vccd1 vccd1 _11905_/B sky130_fd_sc_hd__and3_1
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16424_ input11/X _16424_/D vssd1 vssd1 vccd1 vccd1 _16424_/Q sky130_fd_sc_hd__dfxtp_2
X_13636_ _13636_/A vssd1 vssd1 vccd1 vccd1 _16282_/D sky130_fd_sc_hd__clkbuf_1
X_10848_ _10848_/A vssd1 vssd1 vccd1 vccd1 _15888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13567_ _13561_/C _13562_/C _13564_/Y _13565_/X vssd1 vssd1 vccd1 vccd1 _13568_/C
+ sky130_fd_sc_hd__a211o_1
X_16355_ _16389_/CLK _16355_/D vssd1 vssd1 vccd1 vccd1 _16355_/Q sky130_fd_sc_hd__dfxtp_1
X_10779_ _10779_/A vssd1 vssd1 vccd1 vccd1 _15878_/D sky130_fd_sc_hd__clkbuf_1
X_15306_ _15306_/A vssd1 vssd1 vccd1 vccd1 _15321_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_12518_ _12518_/A _12518_/B vssd1 vssd1 vccd1 vccd1 _12520_/B sky130_fd_sc_hd__nor2_1
X_16286_ _16533_/Q _16286_/D vssd1 vssd1 vccd1 vccd1 _16286_/Q sky130_fd_sc_hd__dfxtp_2
X_13498_ _13498_/A _13498_/B _13503_/A vssd1 vssd1 vccd1 vccd1 _16262_/D sky130_fd_sc_hd__nor3_1
XFILLER_8_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15237_ _15237_/A _15237_/B _15237_/C vssd1 vssd1 vccd1 vccd1 _15238_/C sky130_fd_sc_hd__nand3_1
X_12449_ _16115_/Q _12501_/B _12456_/C vssd1 vssd1 vccd1 vccd1 _12449_/X sky130_fd_sc_hd__and3_1
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15168_ _15169_/B _15169_/C _14954_/X vssd1 vssd1 vccd1 vccd1 _15170_/B sky130_fd_sc_hd__o21ai_1
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _14205_/A _14119_/B _14123_/A vssd1 vssd1 vccd1 vccd1 _16350_/D sky130_fd_sc_hd__nor3_1
XFILLER_125_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07990_ _07991_/B _08204_/A _16571_/Q vssd1 vssd1 vccd1 vccd1 _07992_/A sky130_fd_sc_hd__a21o_1
X_15099_ _15097_/Y _15093_/C _15095_/Y _15096_/X vssd1 vssd1 vccd1 vccd1 _15100_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_113_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09660_ _09529_/X _09656_/B _09659_/Y vssd1 vssd1 vccd1 vccd1 _15667_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ _08730_/A _08611_/B _08621_/B vssd1 vssd1 vccd1 vccd1 _15456_/D sky130_fd_sc_hd__nor3_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09591_ _15657_/Q _09592_/C _09590_/X vssd1 vssd1 vccd1 vccd1 _09591_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08542_ _08542_/A _08542_/B vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__xor2_4
XFILLER_70_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08473_ _08473_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08473_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09025_ _09054_/A _09025_/B _09030_/B vssd1 vssd1 vccd1 vccd1 _15537_/D sky130_fd_sc_hd__nor3_1
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _09925_/X _09927_/B vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__and2b_1
XFILLER_120_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09858_ _15695_/Q _15694_/Q _15693_/Q _09756_/X vssd1 vssd1 vccd1 vccd1 _15705_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08809_ _08809_/A _08809_/B _08809_/C vssd1 vssd1 vccd1 vccd1 _08810_/C sky130_fd_sc_hd__nand3_1
X_09789_ _09744_/X _09787_/B _09788_/Y vssd1 vssd1 vccd1 vccd1 _15693_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11820_ _16026_/Q _11928_/B _11821_/C vssd1 vssd1 vccd1 vccd1 _11820_/X sky130_fd_sc_hd__and3_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11752_/B _11752_/C _11752_/A vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__a21o_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10702_ _15864_/Q _10702_/B _10707_/C vssd1 vssd1 vccd1 vccd1 _10702_/Y sky130_fd_sc_hd__nand3_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _14470_/A vssd1 vssd1 vccd1 vccd1 _16401_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11682_ _11963_/A vssd1 vssd1 vccd1 vccd1 _11805_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13421_ _13705_/A vssd1 vssd1 vccd1 vccd1 _13421_/X sky130_fd_sc_hd__clkbuf_2
X_10633_ _15853_/Q _10679_/B _10639_/C vssd1 vssd1 vccd1 vccd1 _10635_/C sky130_fd_sc_hd__nand3_1
XFILLER_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16140_ _16555_/Q _16140_/D vssd1 vssd1 vccd1 vccd1 _16140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _13349_/Y _13350_/X _13351_/Y _13347_/C vssd1 vssd1 vccd1 vccd1 _13354_/B
+ sky130_fd_sc_hd__o211ai_1
X_10564_ _15839_/Q _10565_/C _10360_/X vssd1 vssd1 vccd1 vccd1 _10566_/A sky130_fd_sc_hd__a21oi_1
X_12303_ _12304_/B _12304_/C _12133_/X vssd1 vssd1 vccd1 vccd1 _12305_/B sky130_fd_sc_hd__o21ai_1
X_16071_ _16118_/CLK _16071_/D vssd1 vssd1 vccd1 vccd1 _16071_/Q sky130_fd_sc_hd__dfxtp_1
X_13283_ _16233_/Q _13336_/B _13283_/C vssd1 vssd1 vccd1 vccd1 _13283_/X sky130_fd_sc_hd__and3_1
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10495_ _10493_/Y _10494_/X _10489_/C _10490_/C vssd1 vssd1 vccd1 vccd1 _10497_/B
+ sky130_fd_sc_hd__o211ai_1
X_15022_ _15023_/B _15023_/C _15023_/A vssd1 vssd1 vccd1 vccd1 _15024_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12234_ _12234_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12236_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12165_ _16075_/Q _12173_/C _12050_/X vssd1 vssd1 vccd1 vccd1 _12165_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11116_ _11152_/C vssd1 vssd1 vccd1 vccd1 _11161_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12096_ _12113_/A _12096_/B _12096_/C vssd1 vssd1 vccd1 vccd1 _12097_/A sky130_fd_sc_hd__and3_1
XFILLER_110_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15924_ _16005_/CLK _15924_/D vssd1 vssd1 vccd1 vccd1 _15924_/Q sky130_fd_sc_hd__dfxtp_1
X_11047_ _11047_/A _11047_/B vssd1 vssd1 vccd1 vccd1 _11048_/B sky130_fd_sc_hd__nor2_1
Xinput9 io_in[8] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_6
X_15855_ _16570_/CLK _15855_/D vssd1 vssd1 vccd1 vccd1 _15855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14806_ _14806_/A vssd1 vssd1 vccd1 vccd1 _15033_/B sky130_fd_sc_hd__clkbuf_2
X_15786_ _15812_/CLK _15786_/D vssd1 vssd1 vccd1 vccd1 _15786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12998_ _13019_/A _12998_/B _12998_/C vssd1 vssd1 vccd1 vccd1 _12999_/A sky130_fd_sc_hd__and3_1
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14737_ _14738_/B _14738_/C _14738_/A vssd1 vssd1 vccd1 vccd1 _14739_/B sky130_fd_sc_hd__a21o_1
X_11949_ _16045_/Q _11950_/C _11726_/X vssd1 vssd1 vccd1 vccd1 _11951_/A sky130_fd_sc_hd__a21oi_1
X_14668_ _14722_/A vssd1 vssd1 vccd1 vccd1 _14707_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16407_ input11/X _16407_/D vssd1 vssd1 vccd1 vccd1 _16407_/Q sky130_fd_sc_hd__dfxtp_2
X_13619_ _13613_/C _13614_/C _13616_/Y _13617_/X vssd1 vssd1 vccd1 vccd1 _13620_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14599_ _14596_/Y _14605_/A _14598_/Y _14594_/C vssd1 vssd1 vccd1 vccd1 _14601_/B
+ sky130_fd_sc_hd__o211a_1
X_16338_ _16346_/CLK _16338_/D vssd1 vssd1 vccd1 vccd1 _16338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16269_ _16533_/Q _16269_/D vssd1 vssd1 vccd1 vccd1 _16269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07973_ _09625_/C _08118_/B vssd1 vssd1 vccd1 vccd1 _07974_/B sky130_fd_sc_hd__xnor2_1
XFILLER_113_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16676__81 vssd1 vssd1 vccd1 vccd1 _16676__81/HI _16752_/A sky130_fd_sc_hd__conb_1
X_09712_ _09717_/C vssd1 vssd1 vccd1 vccd1 _09727_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_101_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09643_ _09643_/A _09643_/B vssd1 vssd1 vccd1 vccd1 _09643_/X sky130_fd_sc_hd__or2_1
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09574_ _09396_/X _09486_/X _09568_/B _09487_/X vssd1 vssd1 vccd1 vccd1 _09575_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _08485_/A _08487_/B _08484_/A vssd1 vssd1 vccd1 vccd1 _08529_/B sky130_fd_sc_hd__a21o_1
XFILLER_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08456_ _08383_/A _08383_/B _08455_/X vssd1 vssd1 vccd1 vccd1 _08497_/B sky130_fd_sc_hd__o21a_2
XFILLER_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08387_ _08388_/A _08388_/B vssd1 vssd1 vccd1 vccd1 _08459_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09008_ _08883_/X _09005_/A _09007_/Y vssd1 vssd1 vccd1 vccd1 _15533_/D sky130_fd_sc_hd__o21a_1
X_10280_ _15804_/Q vssd1 vssd1 vccd1 vccd1 _10285_/B sky130_fd_sc_hd__inv_2
XFILLER_104_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13970_ _13970_/A vssd1 vssd1 vccd1 vccd1 _16329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12921_ _12919_/A _12919_/B _12920_/X vssd1 vssd1 vccd1 vccd1 _16180_/D sky130_fd_sc_hd__a21oi_1
X_15640_ _15812_/CLK _15640_/D vssd1 vssd1 vccd1 vccd1 _15640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _16172_/Q _13022_/B _12852_/C vssd1 vssd1 vccd1 vccd1 _12862_/A sky130_fd_sc_hd__and3_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _16023_/Q _11843_/C _11802_/X vssd1 vssd1 vccd1 vccd1 _11805_/B sky130_fd_sc_hd__a21oi_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _15812_/CLK _15571_/D vssd1 vssd1 vccd1 vccd1 _15571_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _16163_/Q _12792_/C _12619_/X vssd1 vssd1 vccd1 vccd1 _12783_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _11732_/A _11732_/B _11733_/X vssd1 vssd1 vccd1 vccd1 _16012_/D sky130_fd_sc_hd__a21oi_1
X_14522_ _14806_/A vssd1 vssd1 vccd1 vccd1 _14748_/B sky130_fd_sc_hd__buf_2
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11665_ _11663_/Y _11658_/C _11660_/Y _11670_/A vssd1 vssd1 vccd1 vccd1 _11670_/B
+ sky130_fd_sc_hd__a211oi_1
X_14453_ _14454_/B _14454_/C _14454_/A vssd1 vssd1 vccd1 vccd1 _14455_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10616_ _10759_/A _10616_/B vssd1 vssd1 vccd1 vccd1 _10616_/X sky130_fd_sc_hd__or2_1
X_13404_ _13412_/A _13404_/B _13404_/C vssd1 vssd1 vccd1 vccd1 _13405_/A sky130_fd_sc_hd__and3_1
X_14384_ _14437_/A _14389_/C vssd1 vssd1 vccd1 vccd1 _14384_/X sky130_fd_sc_hd__or2_1
X_11596_ _11594_/Y _11589_/C _11592_/Y _11593_/X vssd1 vssd1 vccd1 vccd1 _11597_/C
+ sky130_fd_sc_hd__a211o_1
X_13335_ _16241_/Q _13344_/C _13169_/X vssd1 vssd1 vccd1 vccd1 _13335_/Y sky130_fd_sc_hd__a21oi_1
X_16123_ _16554_/Q _16123_/D vssd1 vssd1 vccd1 vccd1 _16123_/Q sky130_fd_sc_hd__dfxtp_1
X_10547_ _10544_/Y _10546_/X _10541_/C _10542_/C vssd1 vssd1 vccd1 vccd1 _10549_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_115_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16054_ _16118_/CLK _16054_/D vssd1 vssd1 vccd1 vccd1 _16054_/Q sky130_fd_sc_hd__dfxtp_2
X_13266_ _13432_/A _13266_/B _13266_/C vssd1 vssd1 vccd1 vccd1 _13267_/C sky130_fd_sc_hd__or3_1
X_10478_ _15840_/Q vssd1 vssd1 vccd1 vccd1 _10483_/C sky130_fd_sc_hd__inv_2
XFILLER_142_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15005_ _15005_/A _15009_/C vssd1 vssd1 vccd1 vccd1 _15005_/X sky130_fd_sc_hd__or2_1
X_12217_ _16083_/Q _12226_/C _12050_/X vssd1 vssd1 vccd1 vccd1 _12217_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13197_ _13219_/A _13197_/B _13201_/B vssd1 vssd1 vccd1 vccd1 _16219_/D sky130_fd_sc_hd__nor3_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _12148_/A _12148_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12149_/C sky130_fd_sc_hd__nand3_1
XFILLER_110_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12079_ _12100_/C vssd1 vssd1 vccd1 vccd1 _12118_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15907_ _16553_/Q _15907_/D vssd1 vssd1 vccd1 vccd1 _15907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15838_ _16551_/CLK _15838_/D vssd1 vssd1 vccd1 vccd1 _15838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15769_ _15791_/CLK _15769_/D vssd1 vssd1 vccd1 vccd1 _15769_/Q sky130_fd_sc_hd__dfxtp_2
X_08310_ _09278_/A vssd1 vssd1 vccd1 vccd1 _15350_/A sky130_fd_sc_hd__clkbuf_2
X_09290_ _09282_/Y _09288_/X _09289_/Y vssd1 vssd1 vccd1 vccd1 _15593_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _08241_/A _08241_/B vssd1 vssd1 vccd1 vccd1 _08380_/B sky130_fd_sc_hd__xor2_4
XANTENNA_14 _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_25 _10285_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_36 _13443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08172_ _08351_/B _08171_/Y vssd1 vssd1 vccd1 vccd1 _08328_/A sky130_fd_sc_hd__or2b_1
XFILLER_118_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07956_ _16587_/Q _16585_/Q vssd1 vssd1 vccd1 vccd1 _07957_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07887_ _07887_/A _07887_/B vssd1 vssd1 vccd1 vccd1 _07888_/B sky130_fd_sc_hd__nand2_2
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09626_ _09718_/A _09626_/B _09632_/A vssd1 vssd1 vccd1 vccd1 _15661_/D sky130_fd_sc_hd__nor3_1
XFILLER_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09557_ _09557_/A _09557_/B vssd1 vssd1 vccd1 vccd1 _09557_/X sky130_fd_sc_hd__or2_1
XFILLER_102_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08508_ _08509_/A _08509_/B _08509_/C vssd1 vssd1 vccd1 vccd1 _08542_/A sky130_fd_sc_hd__a21oi_4
XFILLER_12_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09488_ _09396_/X _09486_/X _09481_/B _09487_/X vssd1 vssd1 vccd1 vccd1 _09489_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_24_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08439_ _08329_/A _08329_/B _08338_/B vssd1 vssd1 vccd1 vccd1 _08441_/A sky130_fd_sc_hd__a21o_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11450_ _11619_/A vssd1 vssd1 vccd1 vccd1 _11491_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10401_ _15811_/Q _10408_/C _10204_/X vssd1 vssd1 vccd1 vccd1 _10401_/Y sky130_fd_sc_hd__a21oi_1
X_11381_ _15965_/Q _11381_/B _11381_/C vssd1 vssd1 vccd1 vccd1 _11391_/B sky130_fd_sc_hd__and3_1
X_13120_ _16209_/Q _13292_/B _13120_/C vssd1 vssd1 vccd1 vccd1 _13120_/Y sky130_fd_sc_hd__nand3_1
X_10332_ _15798_/Q _10483_/B _10332_/C vssd1 vssd1 vccd1 vccd1 _10337_/A sky130_fd_sc_hd__and3_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13051_ _13051_/A vssd1 vssd1 vccd1 vccd1 _16199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _10260_/Y _10269_/A _10262_/Y _10258_/C vssd1 vssd1 vccd1 vccd1 _10265_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12002_ _16052_/Q _12173_/B _12002_/C vssd1 vssd1 vccd1 vccd1 _12012_/A sky130_fd_sc_hd__and3_1
XFILLER_105_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10194_ _10194_/A vssd1 vssd1 vccd1 vccd1 _15771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16741_ _16741_/A _07848_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_13953_ _13953_/A _13953_/B _13953_/C vssd1 vssd1 vccd1 vccd1 _13954_/C sky130_fd_sc_hd__nand3_1
XFILLER_47_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _16178_/Q _12904_/B _12910_/C vssd1 vssd1 vccd1 vccd1 _12904_/Y sky130_fd_sc_hd__nand3_1
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13884_ _13918_/A _13884_/B _13884_/C vssd1 vssd1 vccd1 vccd1 _13885_/A sky130_fd_sc_hd__and3_1
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15623_ _15812_/CLK _15623_/D vssd1 vssd1 vccd1 vccd1 _15623_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _16170_/Q _13059_/B _12836_/C vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__and3_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15791_/CLK _15554_/D vssd1 vssd1 vccd1 vccd1 _15554_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12766_/A _12766_/B _12766_/C vssd1 vssd1 vccd1 vccd1 _12767_/C sky130_fd_sc_hd__nand3_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _16408_/Q _14547_/C _14339_/X vssd1 vssd1 vccd1 vccd1 _14507_/B sky130_fd_sc_hd__a21oi_1
X_11717_ _11717_/A _11717_/B _11717_/C vssd1 vssd1 vccd1 vccd1 _11718_/A sky130_fd_sc_hd__and3_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15485_ _16570_/CLK _15485_/D vssd1 vssd1 vccd1 vccd1 _15485_/Q sky130_fd_sc_hd__dfxtp_1
X_12697_ _12695_/A _12695_/B _12696_/X vssd1 vssd1 vccd1 vccd1 _16148_/D sky130_fd_sc_hd__a21oi_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11648_ _16001_/Q _11878_/B _11648_/C vssd1 vssd1 vccd1 vccd1 _11648_/Y sky130_fd_sc_hd__nand3_1
X_14436_ _14436_/A _14436_/B vssd1 vssd1 vccd1 vccd1 _14441_/C sky130_fd_sc_hd__nor2_1
XFILLER_128_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11579_ _15992_/Q _11586_/C _11463_/X vssd1 vssd1 vccd1 vccd1 _11582_/B sky130_fd_sc_hd__a21o_1
X_14367_ _14363_/Y _14364_/X _14366_/Y _14361_/C vssd1 vssd1 vccd1 vccd1 _14369_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_10_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16106_ _16118_/CLK _16106_/D vssd1 vssd1 vccd1 vccd1 _16106_/Q sky130_fd_sc_hd__dfxtp_1
X_13318_ _13319_/B _13319_/C _13264_/X vssd1 vssd1 vccd1 vccd1 _13320_/B sky130_fd_sc_hd__o21ai_1
X_14298_ _14291_/C _14292_/C _14295_/Y _14296_/X vssd1 vssd1 vccd1 vccd1 _14299_/C
+ sky130_fd_sc_hd__a211o_1
X_16037_ _16554_/Q _16037_/D vssd1 vssd1 vccd1 vccd1 _16037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13249_ _16228_/Q _13257_/C _13133_/X vssd1 vssd1 vccd1 vccd1 _13249_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07810_ _07811_/A vssd1 vssd1 vccd1 vccd1 _07810_/Y sky130_fd_sc_hd__inv_2
X_08790_ _08790_/A _08790_/B vssd1 vssd1 vccd1 vccd1 _15486_/D sky130_fd_sc_hd__nor2_1
XFILLER_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16646__51 vssd1 vssd1 vccd1 vccd1 _16646__51/HI _16722_/A sky130_fd_sc_hd__conb_1
XFILLER_97_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09411_ _09412_/B _09412_/C _09412_/A vssd1 vssd1 vccd1 vccd1 _09413_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09342_ _09340_/X _09342_/B vssd1 vssd1 vccd1 vccd1 _09342_/X sky130_fd_sc_hd__and2b_1
XFILLER_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09273_ _10789_/B vssd1 vssd1 vccd1 vccd1 _15255_/B sky130_fd_sc_hd__buf_4
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ _08368_/A _08368_/B vssd1 vssd1 vccd1 vccd1 _08225_/B sky130_fd_sc_hd__xor2_2
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08155_ _13943_/A _07911_/B _07910_/A vssd1 vssd1 vccd1 vccd1 _08157_/B sky130_fd_sc_hd__o21ai_4
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08086_ _15489_/Q _08263_/B vssd1 vssd1 vccd1 vccd1 _08266_/B sky130_fd_sc_hd__xnor2_4
XFILLER_146_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08988_ _09054_/A _08988_/B _08993_/B vssd1 vssd1 vccd1 vccd1 _15528_/D sky130_fd_sc_hd__nor3_1
XFILLER_130_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07939_ _08265_/A _07939_/B _07939_/C vssd1 vssd1 vccd1 vccd1 _07941_/A sky130_fd_sc_hd__and3_1
XFILLER_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10950_ _10985_/C vssd1 vssd1 vccd1 vccd1 _10992_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09609_ _09602_/Y _09603_/X _09606_/B vssd1 vssd1 vccd1 vccd1 _09610_/B sky130_fd_sc_hd__o21a_1
X_10881_ _10881_/A _10881_/B vssd1 vssd1 vccd1 vccd1 _10886_/C sky130_fd_sc_hd__nor2_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12620_ _16139_/Q _12628_/C _12619_/X vssd1 vssd1 vccd1 vccd1 _12620_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12551_ input3/X vssd1 vssd1 vccd1 vccd1 _13682_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11502_ _11502_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11503_/B sky130_fd_sc_hd__nor2_1
X_15270_ _15270_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _15274_/C sky130_fd_sc_hd__nor2_1
X_12482_ _12483_/B _12483_/C _12483_/A vssd1 vssd1 vccd1 vccd1 _12484_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11433_ _12849_/A vssd1 vssd1 vccd1 vccd1 _12567_/A sky130_fd_sc_hd__clkbuf_4
X_14221_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__buf_2
XFILLER_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14152_ _14205_/A _14152_/B _14156_/B vssd1 vssd1 vccd1 vccd1 _16355_/D sky130_fd_sc_hd__nor3_1
X_11364_ _11371_/A _11364_/B _11364_/C vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__and3_1
X_10315_ _10315_/A _10315_/B vssd1 vssd1 vccd1 vccd1 _10318_/B sky130_fd_sc_hd__nor2_1
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13103_ _13219_/A _13103_/B _13107_/A vssd1 vssd1 vccd1 vccd1 _16206_/D sky130_fd_sc_hd__nor3_1
X_14083_ _14083_/A vssd1 vssd1 vccd1 vccd1 _16345_/D sky130_fd_sc_hd__clkbuf_1
X_11295_ _15952_/Q _11465_/B _11301_/C vssd1 vssd1 vccd1 vccd1 _11297_/C sky130_fd_sc_hd__nand3_1
XFILLER_112_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13034_ _13034_/A vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__clkbuf_2
X_10246_ _11360_/A vssd1 vssd1 vccd1 vccd1 _10494_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10177_ _15771_/Q _10214_/C _10176_/X vssd1 vssd1 vccd1 vccd1 _10179_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14985_ _14992_/A _14985_/B _14985_/C vssd1 vssd1 vccd1 vccd1 _14986_/A sky130_fd_sc_hd__and3_1
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16724_ _16724_/A _07849_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
X_13936_ _14777_/A vssd1 vssd1 vccd1 vccd1 _14160_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13867_ _13867_/A vssd1 vssd1 vccd1 vccd1 _16314_/D sky130_fd_sc_hd__clkbuf_1
X_15606_ _16551_/CLK _15606_/D vssd1 vssd1 vccd1 vccd1 _15606_/Q sky130_fd_sc_hd__dfxtp_1
X_12818_ _16167_/Q _12818_/B _12828_/C vssd1 vssd1 vccd1 vccd1 _12823_/A sky130_fd_sc_hd__and3_1
XFILLER_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16586_ _16607_/CLK _16586_/D vssd1 vssd1 vccd1 vccd1 _16586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ _16306_/Q _13800_/C _13570_/X vssd1 vssd1 vccd1 vccd1 _13798_/Y sky130_fd_sc_hd__a21oi_1
X_15537_ _15791_/CLK _15537_/D vssd1 vssd1 vccd1 vccd1 _15537_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12749_/A _12753_/C vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__or2_1
XFILLER_148_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15468_ _16551_/CLK _15468_/D vssd1 vssd1 vccd1 vccd1 _15468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14419_ _16395_/Q _14427_/C _14308_/X vssd1 vssd1 vccd1 vccd1 _14419_/Y sky130_fd_sc_hd__a21oi_1
X_15399_ _16085_/Q _16084_/Q _16083_/Q _15397_/X vssd1 vssd1 vccd1 vccd1 _16581_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09960_ _15730_/Q _10003_/B _09966_/C vssd1 vssd1 vccd1 vccd1 _09962_/B sky130_fd_sc_hd__and3_1
XFILLER_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ _08911_/A _08911_/B vssd1 vssd1 vccd1 vccd1 _08912_/B sky130_fd_sc_hd__nor2_1
X_09891_ _09932_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09891_/Y sky130_fd_sc_hd__nor2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08849_/C vssd1 vssd1 vccd1 vccd1 _08866_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _15487_/Q _08943_/B _08779_/C vssd1 vssd1 vccd1 vccd1 _08781_/A sky130_fd_sc_hd__and3_1
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09325_ _09325_/A _09325_/B _09325_/C vssd1 vssd1 vccd1 vccd1 _09326_/C sky130_fd_sc_hd__nand3_1
XFILLER_43_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09256_ _09256_/A _09256_/B _09261_/A vssd1 vssd1 vccd1 vccd1 _15589_/D sky130_fd_sc_hd__nor3_1
X_08207_ _08207_/A vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__inv_2
XFILLER_138_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09187_ _09180_/C _09181_/C _09183_/Y _09194_/A vssd1 vssd1 vccd1 vccd1 _09194_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08138_ _08138_/A _08340_/B vssd1 vssd1 vccd1 vccd1 _08139_/B sky130_fd_sc_hd__xnor2_2
XFILLER_107_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08069_ _16588_/Q _08069_/B vssd1 vssd1 vccd1 vccd1 _08092_/A sky130_fd_sc_hd__xnor2_2
X_10100_ _15756_/Q _10308_/C _10106_/C vssd1 vssd1 vccd1 vccd1 _10100_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11080_ _11078_/Y _11073_/C _11075_/Y _11076_/X vssd1 vssd1 vccd1 vccd1 _11081_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10031_ _15745_/Q _10038_/C _10729_/B vssd1 vssd1 vccd1 vccd1 _10034_/B sky130_fd_sc_hd__a21o_1
XFILLER_49_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ _16450_/Q _14770_/B _14770_/C vssd1 vssd1 vccd1 vccd1 _14780_/B sky130_fd_sc_hd__and3_1
X_11982_ _11998_/A _11982_/B _11982_/C vssd1 vssd1 vccd1 vccd1 _11983_/A sky130_fd_sc_hd__and3_1
XFILLER_44_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13721_ _13738_/C vssd1 vssd1 vccd1 vccd1 _13745_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10933_ _15901_/Q _10934_/C _10874_/X vssd1 vssd1 vccd1 vccd1 _10935_/A sky130_fd_sc_hd__a21oi_1
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16440_ _16595_/CLK _16440_/D vssd1 vssd1 vccd1 vccd1 _16440_/Q sky130_fd_sc_hd__dfxtp_1
X_10864_ _10864_/A _10864_/B _10864_/C vssd1 vssd1 vccd1 vccd1 _10865_/A sky130_fd_sc_hd__and3_1
X_13652_ _13652_/A vssd1 vssd1 vccd1 vccd1 _14777_/A sky130_fd_sc_hd__buf_2
XFILLER_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12603_ _12625_/A _12603_/B _12603_/C vssd1 vssd1 vccd1 vccd1 _12604_/A sky130_fd_sc_hd__and3_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _16389_/CLK _16371_/D vssd1 vssd1 vccd1 vccd1 _16371_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10795_/A vssd1 vssd1 vccd1 vccd1 _15880_/D sky130_fd_sc_hd__clkbuf_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _13583_/A _13583_/B _13583_/C vssd1 vssd1 vccd1 vccd1 _13584_/A sky130_fd_sc_hd__and3_1
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _15327_/A _15327_/B vssd1 vssd1 vccd1 vccd1 _15322_/Y sky130_fd_sc_hd__xnor2_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12534_ _16127_/Q _12578_/C _12368_/X vssd1 vssd1 vccd1 vccd1 _12536_/B sky130_fd_sc_hd__a21oi_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15253_ _16529_/Q _15261_/C _10797_/B vssd1 vssd1 vccd1 vccd1 _15253_/Y sky130_fd_sc_hd__a21oi_1
X_12465_ _12465_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12470_/C sky130_fd_sc_hd__nor2_1
XFILLER_138_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14204_ _14202_/Y _14197_/C _14199_/Y _14209_/A vssd1 vssd1 vccd1 vccd1 _14209_/B
+ sky130_fd_sc_hd__a211oi_1
X_11416_ _11416_/A vssd1 vssd1 vccd1 vccd1 _15968_/D sky130_fd_sc_hd__clkbuf_1
X_15184_ _15184_/A _15184_/B _15184_/C vssd1 vssd1 vccd1 vccd1 _15185_/C sky130_fd_sc_hd__nand3_1
X_12396_ _12392_/Y _12393_/X _12395_/Y _12390_/C vssd1 vssd1 vccd1 vccd1 _12398_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11347_ _15960_/Q _11465_/B _11353_/C vssd1 vssd1 vccd1 vccd1 _11349_/C sky130_fd_sc_hd__nand3_1
XFILLER_4_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ _16353_/Q _14135_/B _14135_/C vssd1 vssd1 vccd1 vccd1 _14135_/Y sky130_fd_sc_hd__nand3_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ _11278_/A _11278_/B vssd1 vssd1 vccd1 vccd1 _11284_/C sky130_fd_sc_hd__nor2_1
X_14066_ _16344_/Q _14289_/B _14072_/C vssd1 vssd1 vccd1 vccd1 _14068_/C sky130_fd_sc_hd__nand3_1
X_10229_ _15795_/Q vssd1 vssd1 vccd1 vccd1 _10235_/C sky130_fd_sc_hd__inv_2
X_13017_ _13014_/Y _13015_/X _13016_/Y _13012_/C vssd1 vssd1 vccd1 vccd1 _13019_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14968_ _16481_/Q _15129_/B _14974_/C vssd1 vssd1 vccd1 vccd1 _14970_/C sky130_fd_sc_hd__nand3_1
XFILLER_35_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16707_ _16707_/A _07808_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_75_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13919_ _13919_/A vssd1 vssd1 vccd1 vccd1 _16322_/D sky130_fd_sc_hd__clkbuf_1
X_14899_ _15415_/A vssd1 vssd1 vccd1 vccd1 _15378_/A sky130_fd_sc_hd__buf_6
XFILLER_63_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16569_ _16570_/CLK _16569_/D vssd1 vssd1 vccd1 vccd1 _16569_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_148_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09110_ _15560_/Q _09192_/B _09110_/C vssd1 vssd1 vccd1 vccd1 _09111_/B sky130_fd_sc_hd__and3_1
XFILLER_31_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09041_ _09041_/A _09041_/B vssd1 vssd1 vccd1 vccd1 _15540_/D sky130_fd_sc_hd__nor2_1
XFILLER_136_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09943_ _09943_/A vssd1 vssd1 vccd1 vccd1 _09943_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _09872_/Y _09879_/A _09869_/C _09870_/C vssd1 vssd1 vccd1 vccd1 _09876_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08825_ _08825_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _08826_/B sky130_fd_sc_hd__nor2_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08756_ _08661_/X _08754_/A _08755_/Y vssd1 vssd1 vccd1 vccd1 _15479_/D sky130_fd_sc_hd__o21a_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08687_ _08730_/A _08687_/B _08691_/B vssd1 vssd1 vccd1 vccd1 _15465_/D sky130_fd_sc_hd__nor3_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09308_ _09792_/A vssd1 vssd1 vccd1 vccd1 _09308_/X sky130_fd_sc_hd__clkbuf_2
X_10580_ _10593_/C vssd1 vssd1 vccd1 vccd1 _10606_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ _09076_/X _09232_/B _09235_/B _09238_/Y vssd1 vssd1 vccd1 vccd1 _15584_/D
+ sky130_fd_sc_hd__o31a_1
X_12250_ _12287_/C vssd1 vssd1 vccd1 vccd1 _12296_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11201_ _11201_/A vssd1 vssd1 vccd1 vccd1 _15937_/D sky130_fd_sc_hd__clkbuf_1
X_12181_ _12181_/A _12181_/B vssd1 vssd1 vccd1 vccd1 _12182_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11132_ _11132_/A vssd1 vssd1 vccd1 vccd1 _15928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15940_ _15365_/A _15940_/D vssd1 vssd1 vccd1 vccd1 _15940_/Q sky130_fd_sc_hd__dfxtp_1
X_11063_ _15920_/Q _11070_/C _10898_/X vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _10008_/Y _10011_/X _10013_/Y vssd1 vssd1 vccd1 vccd1 _15737_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15871_ _16570_/CLK _15871_/D vssd1 vssd1 vccd1 vccd1 _15871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14822_ _16458_/Q _14831_/C _14821_/X vssd1 vssd1 vccd1 vccd1 _14822_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14753_ _14760_/A _14753_/B _14753_/C vssd1 vssd1 vccd1 vccd1 _14754_/A sky130_fd_sc_hd__and3_1
X_11965_ _11979_/C vssd1 vssd1 vccd1 vccd1 _11987_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13704_ _13784_/A _13704_/B _13711_/B vssd1 vssd1 vccd1 vccd1 _16291_/D sky130_fd_sc_hd__nor3_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _10914_/Y _10910_/C _10912_/Y _10913_/X vssd1 vssd1 vccd1 vccd1 _10917_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14684_ _14685_/B _14685_/C _14685_/A vssd1 vssd1 vccd1 vccd1 _14686_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11896_ _16037_/Q _11897_/C _11726_/X vssd1 vssd1 vccd1 vccd1 _11898_/A sky130_fd_sc_hd__a21oi_1
X_16423_ _16595_/CLK _16423_/D vssd1 vssd1 vccd1 vccd1 _16423_/Q sky130_fd_sc_hd__dfxtp_1
X_13635_ _13635_/A _13635_/B _13635_/C vssd1 vssd1 vccd1 vccd1 _13636_/A sky130_fd_sc_hd__and3_1
X_10847_ _10864_/A _10847_/B _10847_/C vssd1 vssd1 vccd1 vccd1 _10848_/A sky130_fd_sc_hd__and3_1
X_16354_ _16389_/CLK _16354_/D vssd1 vssd1 vccd1 vccd1 _16354_/Q sky130_fd_sc_hd__dfxtp_1
X_13566_ _13564_/Y _13565_/X _13561_/C _13562_/C vssd1 vssd1 vccd1 vccd1 _13568_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ _10801_/A _10778_/B _10778_/C vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__and3_1
X_15305_ _15305_/A vssd1 vssd1 vccd1 vccd1 _16538_/D sky130_fd_sc_hd__clkbuf_1
X_12517_ _12517_/A _12526_/B vssd1 vssd1 vccd1 vccd1 _12520_/A sky130_fd_sc_hd__or2_1
XFILLER_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16285_ _16346_/CLK _16285_/D vssd1 vssd1 vccd1 vccd1 _16285_/Q sky130_fd_sc_hd__dfxtp_1
X_13497_ _16263_/Q _13665_/B _13507_/C vssd1 vssd1 vccd1 vccd1 _13503_/A sky130_fd_sc_hd__and3_1
XFILLER_145_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15236_ _15237_/B _15237_/C _15237_/A vssd1 vssd1 vccd1 vccd1 _15238_/B sky130_fd_sc_hd__a21o_1
X_12448_ _16115_/Q _12456_/C _12337_/X vssd1 vssd1 vccd1 vccd1 _12448_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15167_ _15221_/A vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12379_ _16105_/Q _12387_/C _12323_/X vssd1 vssd1 vccd1 vccd1 _12379_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14118_ _16351_/Q _14227_/B _14127_/C vssd1 vssd1 vccd1 vccd1 _14123_/A sky130_fd_sc_hd__and3_1
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15098_ _15095_/Y _15096_/X _15097_/Y _15093_/C vssd1 vssd1 vccd1 vccd1 _15100_/B
+ sky130_fd_sc_hd__o211ai_1
X_14049_ _14047_/A _14047_/B _14048_/X vssd1 vssd1 vccd1 vccd1 _16340_/D sky130_fd_sc_hd__a21oi_1
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08610_ _08592_/C _08593_/C _08605_/Y _08621_/A vssd1 vssd1 vccd1 vccd1 _08621_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09590_ _10294_/C vssd1 vssd1 vccd1 vccd1 _09590_/X sky130_fd_sc_hd__clkbuf_2
X_08541_ _08541_/A _08541_/B vssd1 vssd1 vccd1 vccd1 _08542_/B sky130_fd_sc_hd__nor2_2
XFILLER_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08472_ _08472_/A _08472_/B vssd1 vssd1 vccd1 vccd1 _08475_/A sky130_fd_sc_hd__xnor2_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09024_ _09018_/C _09019_/C _09021_/Y _09030_/A vssd1 vssd1 vccd1 vccd1 _09030_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_117_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09926_ _15722_/Q _09925_/C _08629_/A vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__a21o_1
XFILLER_120_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09857_ _09855_/X _09853_/B _09856_/Y vssd1 vssd1 vccd1 vccd1 _15704_/D sky130_fd_sc_hd__o21a_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _08809_/B _08809_/C _08809_/A vssd1 vssd1 vccd1 vccd1 _08810_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09788_ _09932_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09788_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _10112_/A vssd1 vssd1 vccd1 vccd1 _08916_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _16016_/Q _11750_/B _11757_/C vssd1 vssd1 vccd1 vccd1 _11752_/C sky130_fd_sc_hd__nand3_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _15865_/Q _10929_/B _10701_/C vssd1 vssd1 vccd1 vccd1 _10709_/A sky130_fd_sc_hd__and3_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11681_/A vssd1 vssd1 vccd1 vccd1 _16005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13498_/A _13420_/B _13426_/B vssd1 vssd1 vccd1 vccd1 _16251_/D sky130_fd_sc_hd__nor3_1
XFILLER_139_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10632_ _15853_/Q _10639_/C _10432_/X vssd1 vssd1 vccd1 vccd1 _10635_/B sky130_fd_sc_hd__a21o_1
X_10563_ _10563_/A _10563_/B _10567_/B vssd1 vssd1 vccd1 vccd1 _15836_/D sky130_fd_sc_hd__nor3_1
X_13351_ _16242_/Q _13467_/B _13358_/C vssd1 vssd1 vccd1 vccd1 _13351_/Y sky130_fd_sc_hd__nand3_1
XFILLER_10_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ _12468_/A vssd1 vssd1 vccd1 vccd1 _12343_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16070_ _16118_/CLK _16070_/D vssd1 vssd1 vccd1 vccd1 _16070_/Q sky130_fd_sc_hd__dfxtp_2
X_13282_ _16233_/Q _13292_/C _13169_/X vssd1 vssd1 vccd1 vccd1 _13282_/Y sky130_fd_sc_hd__a21oi_1
X_10494_ _15827_/Q _10494_/B _10494_/C vssd1 vssd1 vccd1 vccd1 _10494_/X sky130_fd_sc_hd__and3_1
XFILLER_108_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ _16490_/Q _15129_/B _15027_/C vssd1 vssd1 vccd1 vccd1 _15023_/C sky130_fd_sc_hd__nand3_1
X_12233_ _12233_/A _12243_/B vssd1 vssd1 vccd1 vccd1 _12236_/A sky130_fd_sc_hd__or2_1
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ _12164_/A vssd1 vssd1 vccd1 vccd1 _16073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _11137_/C vssd1 vssd1 vccd1 vccd1 _11152_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_150_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12095_ _12089_/C _12090_/C _12092_/Y _12093_/X vssd1 vssd1 vccd1 vccd1 _12096_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11046_ _11046_/A _11053_/B vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__or2_1
X_15923_ _15365_/A _15923_/D vssd1 vssd1 vccd1 vccd1 _15923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15854_ _16570_/CLK _15854_/D vssd1 vssd1 vccd1 vccd1 _15854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14805_ _16456_/Q _14808_/C _14694_/X vssd1 vssd1 vccd1 vccd1 _14805_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_92_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15785_ _15812_/CLK _15785_/D vssd1 vssd1 vccd1 vccd1 _15785_/Q sky130_fd_sc_hd__dfxtp_1
X_12997_ _12997_/A _12997_/B _12997_/C vssd1 vssd1 vccd1 vccd1 _12998_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14736_ _16445_/Q _14853_/B _14742_/C vssd1 vssd1 vccd1 vccd1 _14738_/C sky130_fd_sc_hd__nand3_1
XFILLER_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11948_ _11948_/A _11948_/B _11952_/B vssd1 vssd1 vccd1 vccd1 _16043_/D sky130_fd_sc_hd__nor3_1
XFILLER_33_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14667_ _14665_/A _14665_/B _14666_/X vssd1 vssd1 vccd1 vccd1 _16431_/D sky130_fd_sc_hd__a21oi_1
X_11879_ _11876_/Y _11877_/X _11878_/Y _11872_/C vssd1 vssd1 vccd1 vccd1 _11881_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16406_ _16595_/CLK _16406_/D vssd1 vssd1 vccd1 vccd1 _16406_/Q sky130_fd_sc_hd__dfxtp_1
X_13618_ _13616_/Y _13617_/X _13613_/C _13614_/C vssd1 vssd1 vccd1 vccd1 _13620_/B
+ sky130_fd_sc_hd__o211ai_1
X_14598_ _16421_/Q _14598_/B _14603_/C vssd1 vssd1 vccd1 vccd1 _14598_/Y sky130_fd_sc_hd__nand3_1
X_16337_ _16346_/CLK _16337_/D vssd1 vssd1 vccd1 vccd1 _16337_/Q sky130_fd_sc_hd__dfxtp_1
X_13549_ _13583_/A _13549_/B _13549_/C vssd1 vssd1 vccd1 vccd1 _13550_/A sky130_fd_sc_hd__and3_1
XFILLER_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16268_ _16533_/Q _16268_/D vssd1 vssd1 vccd1 vccd1 _16268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15219_ _15271_/A _15223_/C vssd1 vssd1 vccd1 vccd1 _15219_/X sky130_fd_sc_hd__or2_1
XFILLER_133_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16199_ _16555_/Q _16199_/D vssd1 vssd1 vccd1 vccd1 _16199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07972_ _07972_/A _08146_/A vssd1 vssd1 vccd1 vccd1 _08118_/B sky130_fd_sc_hd__xor2_1
XFILLER_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09711_ _15696_/Q vssd1 vssd1 vccd1 vccd1 _09717_/C sky130_fd_sc_hd__inv_2
XFILLER_113_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09642_ _09642_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09642_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09573_ _09394_/X _09568_/B _09572_/X vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__a21oi_1
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _08564_/A _08524_/B vssd1 vssd1 vccd1 vccd1 _08529_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08455_ _08455_/A _08384_/A vssd1 vssd1 vccd1 vccd1 _08455_/X sky130_fd_sc_hd__or2b_1
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08386_ _08386_/A _08386_/B vssd1 vssd1 vccd1 vccd1 _08388_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09007_ _09006_/X _09005_/A _08927_/X vssd1 vssd1 vccd1 vccd1 _09007_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09909_ _09910_/B _09910_/C _09910_/A vssd1 vssd1 vccd1 vccd1 _09911_/B sky130_fd_sc_hd__a21o_1
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12920_ _13032_/A _12925_/C vssd1 vssd1 vccd1 vccd1 _12920_/X sky130_fd_sc_hd__or2_1
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12851_ _16172_/Q _12860_/C _12850_/X vssd1 vssd1 vccd1 vccd1 _12851_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11802_ _12650_/A vssd1 vssd1 vccd1 vccd1 _11802_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _16551_/CLK _15570_/D vssd1 vssd1 vccd1 vccd1 _15570_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12782_/A vssd1 vssd1 vccd1 vccd1 _16161_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _16411_/Q _14524_/C _14411_/X vssd1 vssd1 vccd1 vccd1 _14521_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11733_ _11901_/A _11737_/C vssd1 vssd1 vccd1 vccd1 _11733_/X sky130_fd_sc_hd__or2_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _16400_/Q _14569_/B _14458_/C vssd1 vssd1 vccd1 vccd1 _14454_/C sky130_fd_sc_hd__nand3_1
X_11664_ _11660_/Y _11670_/A _11663_/Y _11658_/C vssd1 vssd1 vccd1 vccd1 _11666_/B
+ sky130_fd_sc_hd__o211a_1
X_13403_ _13401_/Y _13396_/C _13398_/Y _13400_/X vssd1 vssd1 vccd1 vccd1 _13404_/C
+ sky130_fd_sc_hd__a211o_1
X_10615_ _10615_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10616_/B sky130_fd_sc_hd__nor2_1
X_14383_ _14383_/A _14383_/B vssd1 vssd1 vccd1 vccd1 _14389_/C sky130_fd_sc_hd__nor2_1
X_11595_ _11592_/Y _11593_/X _11594_/Y _11589_/C vssd1 vssd1 vccd1 vccd1 _11597_/B
+ sky130_fd_sc_hd__o211ai_1
X_16122_ _16554_/Q _16122_/D vssd1 vssd1 vccd1 vccd1 _16122_/Q sky130_fd_sc_hd__dfxtp_1
X_13334_ _13334_/A vssd1 vssd1 vccd1 vccd1 _16239_/D sky130_fd_sc_hd__clkbuf_1
X_10546_ _15836_/Q _10735_/B _10546_/C vssd1 vssd1 vccd1 vccd1 _10546_/X sky130_fd_sc_hd__and3_1
XFILLER_127_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16053_ _16554_/Q _16053_/D vssd1 vssd1 vccd1 vccd1 _16053_/Q sky130_fd_sc_hd__dfxtp_1
X_13265_ _13266_/B _13266_/C _13264_/X vssd1 vssd1 vccd1 vccd1 _13267_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10477_ _15812_/Q _15811_/Q _15810_/Q _10476_/X vssd1 vssd1 vccd1 vccd1 _15822_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_142_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ _15004_/A _15004_/B vssd1 vssd1 vccd1 vccd1 _15009_/C sky130_fd_sc_hd__nor2_1
X_12216_ _12216_/A vssd1 vssd1 vccd1 vccd1 _16081_/D sky130_fd_sc_hd__clkbuf_1
X_13196_ _13194_/Y _13190_/C _13192_/Y _13201_/A vssd1 vssd1 vccd1 vccd1 _13201_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_2_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12147_ _12148_/B _12148_/C _12148_/A vssd1 vssd1 vccd1 vccd1 _12149_/B sky130_fd_sc_hd__a21o_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12078_ _12093_/C vssd1 vssd1 vccd1 vccd1 _12100_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15906_ _16553_/Q _15906_/D vssd1 vssd1 vccd1 vccd1 _15906_/Q sky130_fd_sc_hd__dfxtp_1
X_11029_ _11036_/A _11029_/B _11029_/C vssd1 vssd1 vccd1 vccd1 _11030_/A sky130_fd_sc_hd__and3_1
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15837_ _16551_/CLK _15837_/D vssd1 vssd1 vccd1 vccd1 _15837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15768_ _15812_/CLK _15768_/D vssd1 vssd1 vccd1 vccd1 _15768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14719_ _14719_/A _14719_/B vssd1 vssd1 vccd1 vccd1 _14724_/C sky130_fd_sc_hd__nor2_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15699_ _15791_/CLK _15699_/D vssd1 vssd1 vccd1 vccd1 _15699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _14675_/A _08048_/B _08239_/X vssd1 vssd1 vccd1 vccd1 _08241_/B sky130_fd_sc_hd__o21a_2
XFILLER_21_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_15 _11150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_26 _15415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08171_ _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08171_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07955_ _16587_/Q _16585_/Q vssd1 vssd1 vccd1 vccd1 _07957_/A sky130_fd_sc_hd__or2_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07886_ _16616_/Q _16614_/Q vssd1 vssd1 vccd1 vccd1 _07887_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ _15664_/Q _09669_/B _09625_/C vssd1 vssd1 vccd1 vccd1 _09632_/A sky130_fd_sc_hd__and3_1
XFILLER_56_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09556_ _09556_/A _09556_/B vssd1 vssd1 vccd1 vccd1 _09556_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08507_ _08443_/A _08443_/B _08506_/X vssd1 vssd1 vccd1 vccd1 _08509_/C sky130_fd_sc_hd__o21a_2
X_09487_ _10618_/A vssd1 vssd1 vccd1 vccd1 _09487_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08438_ _08366_/A _08366_/B _08437_/X vssd1 vssd1 vccd1 vccd1 _08445_/A sky130_fd_sc_hd__a21bo_1
XFILLER_137_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ _08225_/A _08225_/B _08368_/Y vssd1 vssd1 vccd1 vccd1 _08448_/B sky130_fd_sc_hd__a21o_2
XFILLER_137_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10400_ _10400_/A vssd1 vssd1 vccd1 vccd1 _15808_/D sky130_fd_sc_hd__clkbuf_1
X_11380_ _15965_/Q _11381_/C _11158_/X vssd1 vssd1 vccd1 vccd1 _11382_/A sky130_fd_sc_hd__a21oi_1
XFILLER_109_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10331_ _15798_/Q _10362_/C _10176_/X vssd1 vssd1 vccd1 vccd1 _10333_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _15783_/Q _10458_/B _10267_/C vssd1 vssd1 vccd1 vccd1 _10262_/Y sky130_fd_sc_hd__nand3_1
X_13050_ _13072_/A _13050_/B _13050_/C vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__and3_1
XFILLER_127_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12001_ _16052_/Q _12010_/C _12000_/X vssd1 vssd1 vccd1 vccd1 _12001_/Y sky130_fd_sc_hd__a21oi_1
X_10193_ _10250_/A _10193_/B _10193_/C vssd1 vssd1 vccd1 vccd1 _10194_/A sky130_fd_sc_hd__and3_1
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16740_ _16740_/A _07847_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
XFILLER_120_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13952_ _13953_/B _13953_/C _13953_/A vssd1 vssd1 vccd1 vccd1 _13954_/B sky130_fd_sc_hd__a21o_1
XFILLER_101_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12903_ _16179_/Q _13068_/B _12910_/C vssd1 vssd1 vccd1 vccd1 _12903_/X sky130_fd_sc_hd__and3_1
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13883_ _13997_/A _13883_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13884_/C sky130_fd_sc_hd__or3_1
X_15622_ _15812_/CLK _15622_/D vssd1 vssd1 vccd1 vccd1 _15622_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _13682_/A vssd1 vssd1 vccd1 vccd1 _13059_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15791_/CLK _15553_/D vssd1 vssd1 vccd1 vccd1 _15553_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12766_/B _12766_/C _12766_/A vssd1 vssd1 vccd1 vccd1 _12767_/B sky130_fd_sc_hd__a21o_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14539_/C vssd1 vssd1 vccd1 vccd1 _14547_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11716_ _11714_/Y _11709_/C _11711_/Y _11713_/X vssd1 vssd1 vccd1 vccd1 _11717_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _16570_/CLK _15484_/D vssd1 vssd1 vccd1 vccd1 _15484_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12749_/A _12701_/C vssd1 vssd1 vccd1 vccd1 _12696_/X sky130_fd_sc_hd__or2_1
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14435_ _14435_/A _14435_/B vssd1 vssd1 vccd1 vccd1 _14436_/B sky130_fd_sc_hd__nor2_1
X_11647_ _12777_/A vssd1 vssd1 vccd1 vccd1 _11878_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14366_ _16386_/Q _14591_/B _14373_/C vssd1 vssd1 vccd1 vccd1 _14366_/Y sky130_fd_sc_hd__nand3_1
X_11578_ _11666_/A _11578_/B _11582_/A vssd1 vssd1 vccd1 vccd1 _15990_/D sky130_fd_sc_hd__nor3_1
XFILLER_116_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16105_ _16118_/CLK _16105_/D vssd1 vssd1 vccd1 vccd1 _16105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13317_ _13317_/A vssd1 vssd1 vccd1 vccd1 _13354_/A sky130_fd_sc_hd__clkbuf_2
X_10529_ _15821_/Q _15820_/Q _15819_/Q _10476_/X vssd1 vssd1 vccd1 vccd1 _15831_/D
+ sky130_fd_sc_hd__o31a_1
X_14297_ _14295_/Y _14296_/X _14291_/C _14292_/C vssd1 vssd1 vccd1 vccd1 _14299_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16036_ _16554_/Q _16036_/D vssd1 vssd1 vccd1 vccd1 _16036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13248_ _13377_/A vssd1 vssd1 vccd1 vccd1 _13362_/A sky130_fd_sc_hd__buf_2
XFILLER_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13179_ _13176_/Y _13177_/X _13178_/Y _13174_/C vssd1 vssd1 vccd1 vccd1 _13181_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16661__66 vssd1 vssd1 vccd1 vccd1 _16661__66/HI _16737_/A sky130_fd_sc_hd__conb_1
X_09410_ _15620_/Q _09585_/B _09416_/C vssd1 vssd1 vccd1 vccd1 _09412_/C sky130_fd_sc_hd__nand3_1
X_09341_ _15605_/Q _09340_/C _09117_/A vssd1 vssd1 vccd1 vccd1 _09342_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09272_ _15595_/Q _09286_/C _10750_/B vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__a21oi_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08223_ _12247_/A _08018_/B _08222_/X vssd1 vssd1 vccd1 vccd1 _08368_/B sky130_fd_sc_hd__o21a_1
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08154_ _13603_/A _07923_/B _07922_/A vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__o21ai_1
X_08085_ _15471_/Q _15462_/Q vssd1 vssd1 vccd1 vccd1 _08263_/B sky130_fd_sc_hd__xor2_4
XFILLER_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08987_ _08980_/C _08981_/C _08983_/Y _08993_/A vssd1 vssd1 vccd1 vccd1 _08993_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_69_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07938_ _16593_/Q _16591_/Q vssd1 vssd1 vccd1 vccd1 _07939_/C sky130_fd_sc_hd__xor2_1
XFILLER_56_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07869_ _16496_/Q vssd1 vssd1 vccd1 vccd1 _14960_/A sky130_fd_sc_hd__clkinv_2
X_09608_ _09602_/Y _09606_/X _09607_/Y vssd1 vssd1 vccd1 vccd1 _15656_/D sky130_fd_sc_hd__o21a_1
X_10880_ _10880_/A _10880_/B vssd1 vssd1 vccd1 vccd1 _10881_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ _09550_/C vssd1 vssd1 vccd1 vccd1 _09561_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12550_ _16130_/Q _12554_/C _12440_/X vssd1 vssd1 vccd1 vccd1 _12550_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _11501_/A _11509_/B vssd1 vssd1 vccd1 vccd1 _11503_/A sky130_fd_sc_hd__or2_1
XFILLER_8_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _16120_/Q _12600_/B _12487_/C vssd1 vssd1 vccd1 vccd1 _12483_/C sky130_fd_sc_hd__nand3_1
XFILLER_8_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14220_ _14220_/A vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__buf_2
X_11432_ _11432_/A vssd1 vssd1 vccd1 vccd1 _15970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _14149_/Y _14145_/C _14147_/Y _14156_/A vssd1 vssd1 vccd1 vccd1 _14156_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11363_ _11361_/Y _11356_/C _11358_/Y _11359_/X vssd1 vssd1 vccd1 vccd1 _11364_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13102_ _16207_/Q _13102_/B _13112_/C vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__and3_1
X_10314_ _10314_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10318_/A sky130_fd_sc_hd__or2_1
X_14082_ _14090_/A _14082_/B _14082_/C vssd1 vssd1 vccd1 vccd1 _14083_/A sky130_fd_sc_hd__and3_1
X_11294_ _15952_/Q _11301_/C _11181_/X vssd1 vssd1 vccd1 vccd1 _11297_/B sky130_fd_sc_hd__a21o_1
XFILLER_106_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _13031_/A _13031_/B _13032_/X vssd1 vssd1 vccd1 vccd1 _16196_/D sky130_fd_sc_hd__a21oi_1
XFILLER_106_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10245_ _13060_/A vssd1 vssd1 vccd1 vccd1 _11360_/A sky130_fd_sc_hd__buf_4
XFILLER_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10176_ _11233_/A vssd1 vssd1 vccd1 vccd1 _10176_/X sky130_fd_sc_hd__buf_2
XFILLER_94_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14984_ _14982_/Y _14977_/C _14980_/Y _14981_/X vssd1 vssd1 vccd1 vccd1 _14985_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16723_ _16723_/A _07828_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
X_13935_ _13933_/A _13933_/B _13934_/X vssd1 vssd1 vccd1 vccd1 _16324_/D sky130_fd_sc_hd__a21oi_1
XFILLER_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13866_ _13866_/A _13866_/B _13866_/C vssd1 vssd1 vccd1 vccd1 _13867_/A sky130_fd_sc_hd__and3_1
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15605_ _16551_/CLK _15605_/D vssd1 vssd1 vccd1 vccd1 _15605_/Q sky130_fd_sc_hd__dfxtp_1
X_12817_ _16167_/Q _12860_/C _12650_/X vssd1 vssd1 vccd1 vccd1 _12819_/B sky130_fd_sc_hd__a21oi_1
X_16585_ _16595_/CLK _16585_/D vssd1 vssd1 vccd1 vccd1 _16585_/Q sky130_fd_sc_hd__dfxtp_1
X_13797_ _13797_/A vssd1 vssd1 vccd1 vccd1 _16304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15536_ _15791_/CLK _15536_/D vssd1 vssd1 vccd1 vccd1 _15536_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12748_/A _12748_/B vssd1 vssd1 vccd1 vccd1 _12753_/C sky130_fd_sc_hd__nor2_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15467_ _16551_/CLK _15467_/D vssd1 vssd1 vccd1 vccd1 _15467_/Q sky130_fd_sc_hd__dfxtp_1
X_12679_ _12675_/Y _12676_/X _12678_/Y _12673_/C vssd1 vssd1 vccd1 vccd1 _12681_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14418_ _14418_/A vssd1 vssd1 vccd1 vccd1 _16393_/D sky130_fd_sc_hd__clkbuf_1
X_15398_ _16077_/Q _16076_/Q _16075_/Q _15397_/X vssd1 vssd1 vccd1 vccd1 _16580_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14349_ _14349_/A vssd1 vssd1 vccd1 vccd1 _16383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08910_ _10060_/A vssd1 vssd1 vccd1 vccd1 _09074_/A sky130_fd_sc_hd__buf_2
X_16019_ _16554_/Q _16019_/D vssd1 vssd1 vccd1 vccd1 _16019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09890_ _09931_/A _09890_/B vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__and2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _15488_/Q _15487_/Q _15486_/Q _08667_/X vssd1 vssd1 vccd1 vccd1 _15498_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08772_ _09998_/B vssd1 vssd1 vccd1 vccd1 _08943_/B sky130_fd_sc_hd__clkbuf_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09324_ _09325_/B _09325_/C _09325_/A vssd1 vssd1 vccd1 vccd1 _09326_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09255_ _15592_/Q _09448_/B _09255_/C vssd1 vssd1 vccd1 vccd1 _09261_/A sky130_fd_sc_hd__and3_1
XFILLER_21_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08206_ _11287_/A _07998_/B _07997_/B vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__o21ai_1
X_09186_ _09183_/Y _09194_/A _09180_/C _09181_/C vssd1 vssd1 vccd1 vccd1 _09188_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08137_ _08137_/A _08326_/A vssd1 vssd1 vccd1 vccd1 _08340_/B sky130_fd_sc_hd__xnor2_4
XFILLER_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08068_ _12704_/A _08231_/B vssd1 vssd1 vccd1 vccd1 _08069_/B sky130_fd_sc_hd__xnor2_1
XFILLER_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10030_ _10055_/A _10030_/B _10034_/A vssd1 vssd1 vccd1 vccd1 _15742_/D sky130_fd_sc_hd__nor3_1
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11981_ _11974_/C _11975_/C _11977_/Y _11979_/X vssd1 vssd1 vccd1 vccd1 _11982_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13720_ _16608_/Q vssd1 vssd1 vccd1 vccd1 _13738_/C sky130_fd_sc_hd__clkinv_2
X_10932_ _10954_/A _10932_/B _10936_/B vssd1 vssd1 vccd1 vccd1 _15899_/D sky130_fd_sc_hd__nor3_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13651_ _13649_/A _13649_/B _13650_/X vssd1 vssd1 vccd1 vccd1 _16284_/D sky130_fd_sc_hd__a21oi_1
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10863_ _10861_/Y _10855_/C _10857_/Y _10860_/X vssd1 vssd1 vccd1 vccd1 _10864_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12602_ _12602_/A _12602_/B _12602_/C vssd1 vssd1 vccd1 vccd1 _12603_/C sky130_fd_sc_hd__nand3_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _16389_/CLK _16370_/D vssd1 vssd1 vccd1 vccd1 _16370_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13580_/Y _13576_/C _13578_/Y _13579_/X vssd1 vssd1 vccd1 vccd1 _13583_/C
+ sky130_fd_sc_hd__a211o_1
X_10794_ _10801_/A _10794_/B _10794_/C vssd1 vssd1 vccd1 vccd1 _10795_/A sky130_fd_sc_hd__and3_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _16711_/A _15321_/B vssd1 vssd1 vccd1 vccd1 _15327_/B sky130_fd_sc_hd__nand2_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12569_/C vssd1 vssd1 vccd1 vccd1 _12578_/C sky130_fd_sc_hd__clkbuf_2
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ _15252_/A vssd1 vssd1 vccd1 vccd1 _16527_/D sky130_fd_sc_hd__clkbuf_1
X_12464_ _12464_/A _12464_/B vssd1 vssd1 vccd1 vccd1 _12465_/B sky130_fd_sc_hd__nor2_1
XFILLER_126_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14203_ _14199_/Y _14209_/A _14202_/Y _14197_/C vssd1 vssd1 vccd1 vccd1 _14205_/B
+ sky130_fd_sc_hd__o211a_1
X_11415_ _11431_/A _11415_/B _11415_/C vssd1 vssd1 vccd1 vccd1 _11416_/A sky130_fd_sc_hd__and3_1
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15183_ _15184_/B _15184_/C _15184_/A vssd1 vssd1 vccd1 vccd1 _15185_/B sky130_fd_sc_hd__a21o_1
X_12395_ _16106_/Q _12622_/B _12402_/C vssd1 vssd1 vccd1 vccd1 _12395_/Y sky130_fd_sc_hd__nand3_1
X_14134_ _16354_/Q _14185_/B _14135_/C vssd1 vssd1 vccd1 vccd1 _14134_/X sky130_fd_sc_hd__and3_1
X_11346_ _15960_/Q _11353_/C _11181_/X vssd1 vssd1 vccd1 vccd1 _11349_/B sky130_fd_sc_hd__a21o_1
XFILLER_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14065_ _14911_/A vssd1 vssd1 vccd1 vccd1 _14289_/B sky130_fd_sc_hd__clkbuf_2
X_11277_ _11277_/A _11277_/B vssd1 vssd1 vccd1 vccd1 _11278_/B sky130_fd_sc_hd__nor2_1
XFILLER_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13016_ _16194_/Q _13187_/B _13022_/C vssd1 vssd1 vccd1 vccd1 _13016_/Y sky130_fd_sc_hd__nand3_1
XFILLER_140_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10228_ _15767_/Q _15766_/Q _15765_/Q _10227_/X vssd1 vssd1 vccd1 vccd1 _15777_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__or2_1
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14967_ _16481_/Q _14974_/C _14851_/X vssd1 vssd1 vccd1 vccd1 _14970_/B sky130_fd_sc_hd__a21o_1
XFILLER_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16706_ _16706_/A _07807_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13918_ _13918_/A _13918_/B _13918_/C vssd1 vssd1 vccd1 vccd1 _13919_/A sky130_fd_sc_hd__and3_1
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14898_ _14898_/A vssd1 vssd1 vccd1 vccd1 _16468_/D sky130_fd_sc_hd__clkbuf_1
X_16631__36 vssd1 vssd1 vccd1 vccd1 _16631__36/HI _16697_/A sky130_fd_sc_hd__conb_1
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13849_ _13847_/Y _13848_/X _13844_/C _13845_/C vssd1 vssd1 vccd1 vccd1 _13851_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_63_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16568_ _16570_/CLK _16568_/D vssd1 vssd1 vccd1 vccd1 _16568_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15519_ _15791_/CLK _15519_/D vssd1 vssd1 vccd1 vccd1 _15519_/Q sky130_fd_sc_hd__dfxtp_2
X_16499_ _16607_/CLK _16499_/D vssd1 vssd1 vccd1 vccd1 _16499_/Q sky130_fd_sc_hd__dfxtp_1
X_09040_ _09038_/X _09042_/C _09039_/X vssd1 vssd1 vccd1 vccd1 _09041_/B sky130_fd_sc_hd__o21ai_1
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _09955_/C vssd1 vssd1 vccd1 vccd1 _09966_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09873_ _15711_/Q _09914_/B _09873_/C vssd1 vssd1 vccd1 vccd1 _09879_/A sky130_fd_sc_hd__and3_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _08824_/A _08824_/B vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__nor2_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _08663_/X _08754_/A _08711_/X vssd1 vssd1 vccd1 vccd1 _08755_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _08680_/C _08681_/C _08683_/Y _08691_/A vssd1 vssd1 vccd1 vccd1 _08691_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09307_ _09615_/A vssd1 vssd1 vccd1 vccd1 _09307_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09238_ _10065_/A _09244_/C vssd1 vssd1 vccd1 vccd1 _09238_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09169_ _09087_/X _09167_/A _09168_/Y vssd1 vssd1 vccd1 vccd1 _15569_/D sky130_fd_sc_hd__o21a_1
X_11200_ _11208_/A _11200_/B _11200_/C vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__and3_1
XFILLER_107_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12180_ _12180_/A _12187_/B vssd1 vssd1 vccd1 vccd1 _12182_/A sky130_fd_sc_hd__or2_1
XFILLER_108_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11131_ _11148_/A _11131_/B _11131_/C vssd1 vssd1 vccd1 vccd1 _11132_/A sky130_fd_sc_hd__and3_1
XFILLER_135_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11062_ _11097_/A _11062_/B _11066_/A vssd1 vssd1 vccd1 vccd1 _15918_/D sky130_fd_sc_hd__nor3_1
XFILLER_135_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10013_ _10008_/Y _10011_/X _10012_/X vssd1 vssd1 vccd1 vccd1 _10013_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15870_ _16570_/CLK _15870_/D vssd1 vssd1 vccd1 vccd1 _15870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14821_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14821_/X sky130_fd_sc_hd__buf_2
XFILLER_64_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14752_ _14750_/Y _14745_/C _14747_/Y _14748_/X vssd1 vssd1 vccd1 vccd1 _14753_/C
+ sky130_fd_sc_hd__a211o_1
X_11964_ _11964_/A vssd1 vssd1 vccd1 vccd1 _11979_/C sky130_fd_sc_hd__clkbuf_2
X_13703_ _13701_/Y _13696_/C _13699_/Y _13711_/A vssd1 vssd1 vccd1 vccd1 _13711_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_17_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10915_ _10912_/Y _10913_/X _10914_/Y _10910_/C vssd1 vssd1 vccd1 vccd1 _10917_/B
+ sky130_fd_sc_hd__o211ai_1
X_14683_ _16436_/Q _14853_/B _14689_/C vssd1 vssd1 vccd1 vccd1 _14685_/C sky130_fd_sc_hd__nand3_1
XFILLER_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11895_ _11948_/A _11895_/B _11899_/B vssd1 vssd1 vccd1 vccd1 _16035_/D sky130_fd_sc_hd__nor3_1
XFILLER_60_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16422_ _16595_/CLK _16422_/D vssd1 vssd1 vccd1 vccd1 _16422_/Q sky130_fd_sc_hd__dfxtp_1
X_13634_ _13632_/Y _13628_/C _13630_/Y _13631_/X vssd1 vssd1 vccd1 vccd1 _13635_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10846_ _10838_/C _10839_/C _10841_/Y _10844_/X vssd1 vssd1 vccd1 vccd1 _10847_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16353_ _16389_/CLK _16353_/D vssd1 vssd1 vccd1 vccd1 _16353_/Q sky130_fd_sc_hd__dfxtp_1
X_13565_ _16273_/Q _13617_/B _13565_/C vssd1 vssd1 vccd1 vccd1 _13565_/X sky130_fd_sc_hd__and3_1
XFILLER_9_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ _10777_/A _10777_/B _10777_/C vssd1 vssd1 vccd1 vccd1 _10778_/C sky130_fd_sc_hd__nand3_1
X_15304_ _15304_/A _15304_/B vssd1 vssd1 vccd1 vccd1 _15305_/A sky130_fd_sc_hd__and2_1
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12516_ _16125_/Q _12516_/B _12516_/C vssd1 vssd1 vccd1 vccd1 _12526_/B sky130_fd_sc_hd__and3_1
X_16284_ _16346_/CLK _16284_/D vssd1 vssd1 vccd1 vccd1 _16284_/Q sky130_fd_sc_hd__dfxtp_1
X_13496_ _16263_/Q _13538_/C _13495_/X vssd1 vssd1 vccd1 vccd1 _13498_/B sky130_fd_sc_hd__a21oi_1
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15235_ _16526_/Q _15235_/B _15241_/C vssd1 vssd1 vccd1 vccd1 _15237_/C sky130_fd_sc_hd__nand3_1
X_12447_ _12447_/A vssd1 vssd1 vccd1 vccd1 _16113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15166_ _15164_/A _15164_/B _15165_/X vssd1 vssd1 vccd1 vccd1 _16512_/D sky130_fd_sc_hd__a21oi_1
X_12378_ _12378_/A vssd1 vssd1 vccd1 vccd1 _16103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _16351_/Q _14154_/C _14060_/X vssd1 vssd1 vccd1 vccd1 _14119_/B sky130_fd_sc_hd__a21oi_1
X_11329_ _11329_/A _11336_/B vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__or2_1
X_15097_ _16501_/Q _15149_/B _15103_/C vssd1 vssd1 vccd1 vccd1 _15097_/Y sky130_fd_sc_hd__nand3_1
XFILLER_125_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14048_ _14158_/A _14053_/C vssd1 vssd1 vccd1 vccd1 _14048_/X sky130_fd_sc_hd__or2_1
XFILLER_141_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15999_ _16005_/CLK _15999_/D vssd1 vssd1 vccd1 vccd1 _15999_/Q sky130_fd_sc_hd__dfxtp_1
X_08540_ _08540_/A _08540_/B _08540_/C vssd1 vssd1 vccd1 vccd1 _08541_/B sky130_fd_sc_hd__and3_1
XFILLER_36_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08471_ _08512_/A _08512_/B vssd1 vssd1 vccd1 vccd1 _08472_/B sky130_fd_sc_hd__xor2_4
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09023_ _09021_/Y _09030_/A _09018_/C _09019_/C vssd1 vssd1 vccd1 vccd1 _09025_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09925_ _15722_/Q _09966_/B _09925_/C vssd1 vssd1 vccd1 vccd1 _09925_/X sky130_fd_sc_hd__and3_1
XFILLER_131_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09856_ _09207_/X _09853_/B _09750_/X vssd1 vssd1 vccd1 vccd1 _09856_/Y sky130_fd_sc_hd__a21oi_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _15495_/Q _08807_/B _08807_/C vssd1 vssd1 vccd1 vccd1 _08809_/C sky130_fd_sc_hd__nand3_1
X_09787_ _09931_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09788_/B sky130_fd_sc_hd__and2_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _09278_/A vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_26_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _08678_/C vssd1 vssd1 vccd1 vccd1 _08689_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10700_ _14941_/A vssd1 vssd1 vccd1 vccd1 _10929_/B sky130_fd_sc_hd__buf_2
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11717_/A _11680_/B _11680_/C vssd1 vssd1 vccd1 vccd1 _11681_/A sky130_fd_sc_hd__and3_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10631_ _10676_/A _10631_/B _10635_/A vssd1 vssd1 vccd1 vccd1 _15850_/D sky130_fd_sc_hd__nor3_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13350_ _16243_/Q _13350_/B _13358_/C vssd1 vssd1 vccd1 vccd1 _13350_/X sky130_fd_sc_hd__and3_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10562_ _10560_/Y _10556_/C _10558_/Y _10567_/A vssd1 vssd1 vccd1 vccd1 _10567_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _12299_/A _12299_/B _12300_/X vssd1 vssd1 vccd1 vccd1 _16092_/D sky130_fd_sc_hd__a21oi_1
XFILLER_139_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13281_ _13281_/A vssd1 vssd1 vccd1 vccd1 _16231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10493_ _15827_/Q _10494_/C _10492_/X vssd1 vssd1 vccd1 vccd1 _10493_/Y sky130_fd_sc_hd__a21oi_1
X_15020_ _16490_/Q _15027_/C _14851_/X vssd1 vssd1 vccd1 vccd1 _15023_/B sky130_fd_sc_hd__a21o_1
X_12232_ _16085_/Q _12232_/B _12232_/C vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__and3_1
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _12170_/A _12163_/B _12163_/C vssd1 vssd1 vccd1 vccd1 _12164_/A sky130_fd_sc_hd__and3_1
XFILLER_123_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11114_ _11128_/C vssd1 vssd1 vccd1 vccd1 _11137_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12094_ _12092_/Y _12093_/X _12089_/C _12090_/C vssd1 vssd1 vccd1 vccd1 _12096_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11045_ _15917_/Q _11099_/B _11045_/C vssd1 vssd1 vccd1 vccd1 _11053_/B sky130_fd_sc_hd__and3_1
X_15922_ _16005_/CLK _15922_/D vssd1 vssd1 vccd1 vccd1 _15922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15853_ _16570_/CLK _15853_/D vssd1 vssd1 vccd1 vccd1 _15853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14804_ _14804_/A vssd1 vssd1 vccd1 vccd1 _16454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15784_ _15812_/CLK _15784_/D vssd1 vssd1 vccd1 vccd1 _15784_/Q sky130_fd_sc_hd__dfxtp_1
X_12996_ _12997_/B _12997_/C _12997_/A vssd1 vssd1 vccd1 vccd1 _12998_/B sky130_fd_sc_hd__a21o_1
XFILLER_92_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11947_ _11945_/Y _11940_/C _11942_/Y _11952_/A vssd1 vssd1 vccd1 vccd1 _11952_/B
+ sky130_fd_sc_hd__a211oi_1
X_14735_ _16445_/Q _14742_/C _14567_/X vssd1 vssd1 vccd1 vccd1 _14738_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14666_ _14720_/A _14671_/C vssd1 vssd1 vccd1 vccd1 _14666_/X sky130_fd_sc_hd__or2_1
X_11878_ _16033_/Q _11878_/B _11878_/C vssd1 vssd1 vccd1 vccd1 _11878_/Y sky130_fd_sc_hd__nand3_1
X_13617_ _16281_/Q _13617_/B _13617_/C vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__and3_1
X_16405_ _16607_/CLK _16405_/D vssd1 vssd1 vccd1 vccd1 _16405_/Q sky130_fd_sc_hd__dfxtp_1
X_10829_ _10844_/C vssd1 vssd1 vccd1 vccd1 _10852_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14597_ _16422_/Q _14710_/B _14597_/C vssd1 vssd1 vccd1 vccd1 _14605_/A sky130_fd_sc_hd__and3_1
XFILLER_41_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13548_ _13717_/A _13548_/B _13548_/C vssd1 vssd1 vccd1 vccd1 _13549_/C sky130_fd_sc_hd__or3_1
X_16336_ _16389_/CLK _16336_/D vssd1 vssd1 vccd1 vccd1 _16336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16267_ _16533_/Q _16267_/D vssd1 vssd1 vccd1 vccd1 _16267_/Q sky130_fd_sc_hd__dfxtp_1
X_13479_ _16261_/Q _13645_/B _13479_/C vssd1 vssd1 vccd1 vccd1 _13488_/B sky130_fd_sc_hd__and3_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15218_ _15218_/A _15218_/B vssd1 vssd1 vccd1 vccd1 _15223_/C sky130_fd_sc_hd__nor2_1
X_16198_ _16555_/Q _16198_/D vssd1 vssd1 vccd1 vccd1 _16198_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _16510_/Q _15149_/B _15155_/C vssd1 vssd1 vccd1 vccd1 _15149_/Y sky130_fd_sc_hd__nand3_1
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07971_ _09802_/C _08147_/B vssd1 vssd1 vccd1 vccd1 _08146_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09710_ _15668_/Q _15667_/Q _15666_/Q _09536_/X vssd1 vssd1 vccd1 vccd1 _15678_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09641_ _15667_/Q _09641_/B _09648_/C vssd1 vssd1 vccd1 vccd1 _09643_/B sky130_fd_sc_hd__and3_1
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09572_ _10418_/A vssd1 vssd1 vccd1 vccd1 _09572_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08523_ _15451_/Q _08561_/B _15307_/C vssd1 vssd1 vccd1 vccd1 _08524_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08454_ _08454_/A _08454_/B _08373_/B vssd1 vssd1 vccd1 vccd1 _08497_/A sky130_fd_sc_hd__or3b_1
XFILLER_35_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08385_ _16534_/Q _16532_/Q _08385_/C vssd1 vssd1 vccd1 vccd1 _08388_/A sky130_fd_sc_hd__and3_1
XFILLER_136_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09006_ _09207_/A vssd1 vssd1 vccd1 vccd1 _09006_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16667__72 vssd1 vssd1 vccd1 vccd1 _16667__72/HI _16743_/A sky130_fd_sc_hd__conb_1
X_09908_ _15719_/Q _09992_/B _09914_/C vssd1 vssd1 vccd1 vccd1 _09910_/C sky130_fd_sc_hd__nand3_1
XFILLER_86_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09839_ _09835_/Y _09847_/A _09838_/Y _09831_/C vssd1 vssd1 vccd1 vccd1 _09841_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ _13979_/A vssd1 vssd1 vccd1 vccd1 _12850_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11801_ _11836_/C vssd1 vssd1 vccd1 vccd1 _11843_/C sky130_fd_sc_hd__clkbuf_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12781_ _12788_/A _12781_/B _12781_/C vssd1 vssd1 vccd1 vccd1 _12782_/A sky130_fd_sc_hd__and3_1
XFILLER_42_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14520_/A vssd1 vssd1 vccd1 vccd1 _16409_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11732_ _11732_/A _11732_/B vssd1 vssd1 vccd1 vccd1 _11737_/C sky130_fd_sc_hd__nor2_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _16400_/Q _14458_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14454_/B sky130_fd_sc_hd__a21o_1
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11663_ _16003_/Q _11780_/B _11668_/C vssd1 vssd1 vccd1 vccd1 _11663_/Y sky130_fd_sc_hd__nand3_1
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13398_/Y _13400_/X _13401_/Y _13396_/C vssd1 vssd1 vccd1 vccd1 _13404_/B
+ sky130_fd_sc_hd__o211ai_1
X_10614_ _10614_/A _10614_/B vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__nor2_1
X_14382_ _14382_/A _14382_/B vssd1 vssd1 vccd1 vccd1 _14383_/B sky130_fd_sc_hd__nor2_1
X_11594_ _15993_/Q _11594_/B _11594_/C vssd1 vssd1 vccd1 vccd1 _11594_/Y sky130_fd_sc_hd__nand3_1
X_16121_ _16554_/Q _16121_/D vssd1 vssd1 vccd1 vccd1 _16121_/Q sky130_fd_sc_hd__dfxtp_1
X_13333_ _13354_/A _13333_/B _13333_/C vssd1 vssd1 vccd1 vccd1 _13334_/A sky130_fd_sc_hd__and3_1
XFILLER_127_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10545_ _11360_/A vssd1 vssd1 vccd1 vccd1 _10735_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16052_ _16554_/Q _16052_/D vssd1 vssd1 vccd1 vccd1 _16052_/Q sky130_fd_sc_hd__dfxtp_1
X_13264_ _13264_/A vssd1 vssd1 vccd1 vccd1 _13264_/X sky130_fd_sc_hd__clkbuf_2
X_10476_ _14615_/A vssd1 vssd1 vccd1 vccd1 _10476_/X sky130_fd_sc_hd__clkbuf_2
X_15003_ _15003_/A _15003_/B vssd1 vssd1 vccd1 vccd1 _15004_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12215_ _12222_/A _12215_/B _12215_/C vssd1 vssd1 vccd1 vccd1 _12216_/A sky130_fd_sc_hd__and3_1
X_13195_ _13192_/Y _13201_/A _13194_/Y _13190_/C vssd1 vssd1 vccd1 vccd1 _13197_/B
+ sky130_fd_sc_hd__o211a_1
X_12146_ _16072_/Q _12318_/B _12152_/C vssd1 vssd1 vccd1 vccd1 _12148_/C sky130_fd_sc_hd__nand3_1
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12077_ _16579_/Q vssd1 vssd1 vccd1 vccd1 _12093_/C sky130_fd_sc_hd__clkinv_2
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11028_ _11026_/Y _11021_/C _11024_/Y _11025_/X vssd1 vssd1 vccd1 vccd1 _11029_/C
+ sky130_fd_sc_hd__a211o_1
X_15905_ _16553_/Q _15905_/D vssd1 vssd1 vccd1 vccd1 _15905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15836_ _16570_/CLK _15836_/D vssd1 vssd1 vccd1 vccd1 _15836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15767_ _15812_/CLK _15767_/D vssd1 vssd1 vccd1 vccd1 _15767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12979_ _13032_/A _12984_/C vssd1 vssd1 vccd1 vccd1 _12979_/X sky130_fd_sc_hd__or2_1
XFILLER_45_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14718_ _14718_/A _14718_/B vssd1 vssd1 vccd1 vccd1 _14719_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15698_ _15791_/CLK _15698_/D vssd1 vssd1 vccd1 vccd1 _15698_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ _14645_/Y _14646_/X _14648_/Y _14643_/C vssd1 vssd1 vccd1 vccd1 _14651_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_16 _11233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16319_ _16346_/CLK _16319_/D vssd1 vssd1 vccd1 vccd1 _16319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07954_ _16589_/Q vssd1 vssd1 vccd1 vccd1 _12646_/A sky130_fd_sc_hd__clkinv_2
X_07885_ _16616_/Q _16614_/Q vssd1 vssd1 vccd1 vccd1 _07887_/A sky130_fd_sc_hd__or2_1
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09624_ _15664_/Q _09648_/C _09493_/X vssd1 vssd1 vccd1 vccd1 _09626_/B sky130_fd_sc_hd__a21oi_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09555_ _15649_/Q _09641_/B _09561_/C vssd1 vssd1 vccd1 vccd1 _09557_/B sky130_fd_sc_hd__and3_1
XFILLER_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08506_ _08441_/A _08441_/B _08444_/B vssd1 vssd1 vccd1 vccd1 _08506_/X sky130_fd_sc_hd__a21o_1
X_09486_ _09792_/A vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08437_ _08437_/A _08367_/A vssd1 vssd1 vccd1 vccd1 _08437_/X sky130_fd_sc_hd__or2b_1
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08368_ _08368_/A _08368_/B vssd1 vssd1 vccd1 vccd1 _08368_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08299_ _08299_/A _08298_/A vssd1 vssd1 vccd1 vccd1 _08300_/B sky130_fd_sc_hd__or2b_1
XFILLER_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10330_ _10355_/C vssd1 vssd1 vccd1 vccd1 _10362_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_124_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10261_ _15784_/Q _10402_/B _10261_/C vssd1 vssd1 vccd1 vccd1 _10269_/A sky130_fd_sc_hd__and3_1
X_12000_ _12567_/A vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10192_ _10186_/C _10187_/C _10189_/Y _10190_/X vssd1 vssd1 vccd1 vccd1 _10193_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13951_ _16328_/Q _14010_/B _13958_/C vssd1 vssd1 vccd1 vccd1 _13953_/C sky130_fd_sc_hd__nand3_1
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12902_ _16179_/Q _12910_/C _12901_/X vssd1 vssd1 vccd1 vccd1 _12902_/Y sky130_fd_sc_hd__a21oi_1
X_13882_ _13883_/B _13883_/C _13829_/X vssd1 vssd1 vccd1 vccd1 _13884_/B sky130_fd_sc_hd__o21ai_1
XFILLER_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15621_ _15812_/CLK _15621_/D vssd1 vssd1 vccd1 vccd1 _15621_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ _16170_/Q _12836_/C _12723_/X vssd1 vssd1 vccd1 vccd1 _12833_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _16160_/Q _12881_/B _12770_/C vssd1 vssd1 vccd1 vccd1 _12766_/C sky130_fd_sc_hd__nand3_1
X_15552_ _16551_/CLK _15552_/D vssd1 vssd1 vccd1 vccd1 _15552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11715_ _11711_/Y _11713_/X _11714_/Y _11709_/C vssd1 vssd1 vccd1 vccd1 _11717_/B
+ sky130_fd_sc_hd__o211ai_1
X_14503_ _14524_/C vssd1 vssd1 vccd1 vccd1 _14539_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15483_ _16570_/CLK _15483_/D vssd1 vssd1 vccd1 vccd1 _15483_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12695_/A _12695_/B vssd1 vssd1 vccd1 vccd1 _12701_/C sky130_fd_sc_hd__nor2_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11646_ _15241_/B vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__buf_4
X_14434_ _14434_/A _14441_/B vssd1 vssd1 vccd1 vccd1 _14436_/A sky130_fd_sc_hd__or2_1
XFILLER_128_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14365_ _14647_/A vssd1 vssd1 vccd1 vccd1 _14591_/B sky130_fd_sc_hd__clkbuf_2
X_11577_ _15991_/Q _11688_/B _11586_/C vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__and3_1
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16104_ _16118_/CLK _16104_/D vssd1 vssd1 vccd1 vccd1 _16104_/Q sky130_fd_sc_hd__dfxtp_1
X_13316_ _13314_/A _13314_/B _13315_/X vssd1 vssd1 vccd1 vccd1 _16236_/D sky130_fd_sc_hd__a21oi_1
X_10528_ _10526_/X _10524_/B _10527_/Y vssd1 vssd1 vccd1 vccd1 _15830_/D sky130_fd_sc_hd__o21a_1
X_14296_ _16377_/Q _14458_/B _14296_/C vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__and3_1
X_16035_ _16118_/CLK _16035_/D vssd1 vssd1 vccd1 vccd1 _16035_/Q sky130_fd_sc_hd__dfxtp_1
X_13247_ _13247_/A vssd1 vssd1 vccd1 vccd1 _16226_/D sky130_fd_sc_hd__clkbuf_1
X_10459_ _10455_/Y _10465_/A _10458_/Y _10451_/C vssd1 vssd1 vccd1 vccd1 _10461_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ _16217_/Q _13292_/B _13178_/C vssd1 vssd1 vccd1 vccd1 _13178_/Y sky130_fd_sc_hd__nand3_1
X_12129_ _12183_/A _12135_/C vssd1 vssd1 vccd1 vccd1 _12129_/X sky130_fd_sc_hd__or2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15819_ _16551_/CLK _15819_/D vssd1 vssd1 vccd1 vccd1 _15819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09340_ _15605_/Q _09472_/B _09340_/C vssd1 vssd1 vccd1 vccd1 _09340_/X sky130_fd_sc_hd__and3_1
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09271_ _09271_/A vssd1 vssd1 vccd1 vccd1 _10750_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08222_ _12364_/A _08222_/B vssd1 vssd1 vccd1 vccd1 _08222_/X sky130_fd_sc_hd__or2_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08153_ _13435_/A _07930_/B _07933_/A vssd1 vssd1 vccd1 vccd1 _08330_/A sky130_fd_sc_hd__o21bai_1
XFILLER_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08084_ _16523_/Q vssd1 vssd1 vccd1 vccd1 _15121_/A sky130_fd_sc_hd__clkinv_2
XFILLER_130_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _08983_/Y _08993_/A _08980_/C _08981_/C vssd1 vssd1 vccd1 vccd1 _08988_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16637__42 vssd1 vssd1 vccd1 vccd1 _16637__42/HI _16713_/A sky130_fd_sc_hd__conb_1
XFILLER_69_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07937_ _16534_/Q _16532_/Q vssd1 vssd1 vccd1 vccd1 _07939_/B sky130_fd_sc_hd__or2_2
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07868_ _16595_/Q vssd1 vssd1 vccd1 vccd1 _12987_/A sky130_fd_sc_hd__clkinv_2
XFILLER_113_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09607_ _09602_/Y _09606_/X _09530_/X vssd1 vssd1 vccd1 vccd1 _09607_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07799_ _07799_/A vssd1 vssd1 vccd1 vccd1 _07799_/Y sky130_fd_sc_hd__inv_2
X_09538_ _09541_/C vssd1 vssd1 vccd1 vccd1 _09550_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _09468_/X _09467_/Y _09424_/X vssd1 vssd1 vccd1 vccd1 _09469_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ _15981_/Q _11668_/B _11500_/C vssd1 vssd1 vccd1 vccd1 _11509_/B sky130_fd_sc_hd__and3_1
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12480_ _16120_/Q _12487_/C _12316_/X vssd1 vssd1 vccd1 vccd1 _12483_/B sky130_fd_sc_hd__a21o_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11431_ _11431_/A _11431_/B _11431_/C vssd1 vssd1 vccd1 vccd1 _11432_/A sky130_fd_sc_hd__and3_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14150_ _14147_/Y _14156_/A _14149_/Y _14145_/C vssd1 vssd1 vccd1 vccd1 _14152_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ _11358_/Y _11359_/X _11361_/Y _11356_/C vssd1 vssd1 vccd1 vccd1 _11364_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_125_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13101_ _16207_/Q _13143_/C _12933_/X vssd1 vssd1 vccd1 vccd1 _13103_/B sky130_fd_sc_hd__a21oi_1
X_10313_ _15794_/Q _10313_/B _10313_/C vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__and3_1
XFILLER_98_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14081_ _14079_/Y _14075_/C _14077_/Y _14078_/X vssd1 vssd1 vccd1 vccd1 _14082_/C
+ sky130_fd_sc_hd__a211o_1
X_11293_ _11379_/A _11293_/B _11297_/A vssd1 vssd1 vccd1 vccd1 _15950_/D sky130_fd_sc_hd__nor3_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13032_ _13032_/A _13036_/C vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__or2_1
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10244_ _15782_/Q _10247_/C _10243_/X vssd1 vssd1 vccd1 vccd1 _10244_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10175_ _12932_/A vssd1 vssd1 vccd1 vccd1 _11233_/A sky130_fd_sc_hd__buf_4
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14983_ _14980_/Y _14981_/X _14982_/Y _14977_/C vssd1 vssd1 vccd1 vccd1 _14985_/B
+ sky130_fd_sc_hd__o211ai_1
X_16722_ _16722_/A _07827_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
X_13934_ _14158_/A _13939_/C vssd1 vssd1 vccd1 vccd1 _13934_/X sky130_fd_sc_hd__or2_1
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13865_ _13863_/Y _13859_/C _13861_/Y _13862_/X vssd1 vssd1 vccd1 vccd1 _13866_/C
+ sky130_fd_sc_hd__a211o_1
X_15604_ _16551_/CLK _15604_/D vssd1 vssd1 vccd1 vccd1 _15604_/Q sky130_fd_sc_hd__dfxtp_1
X_12816_ _12852_/C vssd1 vssd1 vccd1 vccd1 _12860_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16584_ _16595_/CLK _16584_/D vssd1 vssd1 vccd1 vccd1 _16584_/Q sky130_fd_sc_hd__dfxtp_1
X_13796_ _13811_/A _13796_/B _13796_/C vssd1 vssd1 vccd1 vccd1 _13797_/A sky130_fd_sc_hd__and3_1
X_15535_ _15791_/CLK _15535_/D vssd1 vssd1 vccd1 vccd1 _15535_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12747_/A _12747_/B vssd1 vssd1 vccd1 vccd1 _12748_/B sky130_fd_sc_hd__nor2_1
XFILLER_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _16146_/Q _12904_/B _12685_/C vssd1 vssd1 vccd1 vccd1 _12678_/Y sky130_fd_sc_hd__nand3_1
X_15466_ _16551_/CLK _15466_/D vssd1 vssd1 vccd1 vccd1 _15466_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11629_ _15999_/Q _11688_/B _11638_/C vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__and3_1
X_14417_ _14424_/A _14417_/B _14417_/C vssd1 vssd1 vccd1 vccd1 _14418_/A sky130_fd_sc_hd__and3_1
XFILLER_128_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15397_ _15409_/A vssd1 vssd1 vccd1 vccd1 _15397_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14348_ _14369_/A _14348_/B _14348_/C vssd1 vssd1 vccd1 vccd1 _14349_/A sky130_fd_sc_hd__and3_1
XFILLER_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14279_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14296_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16018_ _16554_/Q _16018_/D vssd1 vssd1 vccd1 vccd1 _16018_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08661_/X _08838_/A _08839_/Y vssd1 vssd1 vccd1 vccd1 _15497_/D sky130_fd_sc_hd__o21a_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _15487_/Q _08779_/C _08604_/X vssd1 vssd1 vccd1 vccd1 _08771_/Y sky130_fd_sc_hd__a21oi_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09323_ _15602_/Q _09364_/B _09329_/C vssd1 vssd1 vccd1 vccd1 _09325_/C sky130_fd_sc_hd__nand3_1
XFILLER_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09254_ _09801_/A vssd1 vssd1 vccd1 vccd1 _09448_/B sky130_fd_sc_hd__buf_2
XFILLER_138_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08205_ _08357_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ _15577_/Q _15341_/B _09192_/C vssd1 vssd1 vccd1 vccd1 _09194_/A sky130_fd_sc_hd__and3_1
XFILLER_119_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08136_ _08136_/A _08325_/A vssd1 vssd1 vccd1 vccd1 _08326_/A sky130_fd_sc_hd__xor2_4
XFILLER_135_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08067_ _08245_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08231_/B sky130_fd_sc_hd__xor2_4
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08969_ _10697_/A vssd1 vssd1 vccd1 vccd1 _09400_/A sky130_fd_sc_hd__buf_2
XFILLER_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11980_ _11977_/Y _11979_/X _11974_/C _11975_/C vssd1 vssd1 vccd1 vccd1 _11982_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_72_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ _10929_/Y _10925_/C _10927_/Y _10936_/A vssd1 vssd1 vccd1 vccd1 _10936_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10862_ _10857_/Y _10860_/X _10861_/Y _10855_/C vssd1 vssd1 vccd1 vccd1 _10864_/B
+ sky130_fd_sc_hd__o211ai_1
X_13650_ _13879_/A _13656_/C vssd1 vssd1 vccd1 vccd1 _13650_/X sky130_fd_sc_hd__or2_1
XFILLER_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12602_/B _12602_/C _12602_/A vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__a21o_1
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _13578_/Y _13579_/X _13580_/Y _13576_/C vssd1 vssd1 vccd1 vccd1 _13583_/B
+ sky130_fd_sc_hd__o211ai_1
X_10793_ _10791_/Y _10785_/C _10788_/Y _10789_/X vssd1 vssd1 vccd1 vccd1 _10794_/C
+ sky130_fd_sc_hd__a211o_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _12554_/C vssd1 vssd1 vccd1 vccd1 _12569_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15320_ _15320_/A vssd1 vssd1 vccd1 vccd1 _15320_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15251_ _15258_/A _15251_/B _15251_/C vssd1 vssd1 vccd1 vccd1 _15252_/A sky130_fd_sc_hd__and3_1
X_12463_ _12463_/A _12470_/B vssd1 vssd1 vccd1 vccd1 _12465_/A sky130_fd_sc_hd__or2_1
XFILLER_138_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11414_ _11407_/C _11408_/C _11410_/Y _11412_/X vssd1 vssd1 vccd1 vccd1 _11415_/C
+ sky130_fd_sc_hd__a211o_1
X_14202_ _16363_/Q _14318_/B _14207_/C vssd1 vssd1 vccd1 vccd1 _14202_/Y sky130_fd_sc_hd__nand3_1
X_15182_ _16517_/Q _15235_/B _15188_/C vssd1 vssd1 vccd1 vccd1 _15184_/C sky130_fd_sc_hd__nand3_1
X_12394_ _13242_/A vssd1 vssd1 vccd1 vccd1 _12622_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_125_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14133_ _16354_/Q _14135_/C _14132_/X vssd1 vssd1 vccd1 vccd1 _14133_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11345_ _11379_/A _11345_/B _11349_/A vssd1 vssd1 vccd1 vccd1 _15958_/D sky130_fd_sc_hd__nor3_1
XFILLER_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14064_ _16344_/Q _14072_/C _14008_/X vssd1 vssd1 vccd1 vccd1 _14068_/B sky130_fd_sc_hd__a21o_1
X_11276_ _11276_/A _11284_/B vssd1 vssd1 vccd1 vccd1 _11278_/A sky130_fd_sc_hd__or2_1
XFILLER_140_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13015_ _16195_/Q _13068_/B _13022_/C vssd1 vssd1 vccd1 vccd1 _13015_/X sky130_fd_sc_hd__and3_1
X_10227_ _14615_/A vssd1 vssd1 vccd1 vccd1 _10227_/X sky130_fd_sc_hd__buf_2
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10158_ _15767_/Q _10313_/C _10158_/C vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__and3_1
XFILLER_67_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10089_ _10145_/A _10089_/B _10089_/C vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__and3_1
X_14966_ _15053_/A _14966_/B _14970_/A vssd1 vssd1 vccd1 vccd1 _16479_/D sky130_fd_sc_hd__nor3_1
XFILLER_48_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ _16705_/A _07805_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13917_ _13915_/Y _13911_/C _13913_/Y _13914_/X vssd1 vssd1 vccd1 vccd1 _13918_/C
+ sky130_fd_sc_hd__a211o_1
X_14897_ _14936_/A _14897_/B _14897_/C vssd1 vssd1 vccd1 vccd1 _14898_/A sky130_fd_sc_hd__and3_1
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13848_ _16313_/Q _13900_/B _13848_/C vssd1 vssd1 vccd1 vccd1 _13848_/X sky130_fd_sc_hd__and3_1
XFILLER_16_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16567_ _16570_/CLK _16567_/D vssd1 vssd1 vccd1 vccd1 _16567_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13779_ _13800_/C vssd1 vssd1 vccd1 vccd1 _13815_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15518_ _15791_/CLK _15518_/D vssd1 vssd1 vccd1 vccd1 _15518_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16498_ _16607_/CLK _16498_/D vssd1 vssd1 vccd1 vccd1 _16498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15449_ _16570_/CLK _15449_/D vssd1 vssd1 vccd1 vccd1 _15449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09941_ _09945_/C vssd1 vssd1 vccd1 vccd1 _09955_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _15711_/Q _09873_/C _08604_/A vssd1 vssd1 vccd1 vccd1 _09872_/Y sky130_fd_sc_hd__a21oi_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08823_/A _08823_/B vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__or2_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08754_ _08754_/A _08754_/B vssd1 vssd1 vccd1 vccd1 _15478_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _08683_/Y _08691_/A _08680_/C _08681_/C vssd1 vssd1 vccd1 vccd1 _08687_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09306_ _09299_/X _09296_/B _09305_/Y vssd1 vssd1 vccd1 vccd1 _15595_/D sky130_fd_sc_hd__o21a_1
XFILLER_22_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09237_ _09232_/B _09235_/B _09117_/X vssd1 vssd1 vccd1 vccd1 _09244_/C sky130_fd_sc_hd__o21a_1
X_09168_ _09006_/X _09167_/A _09129_/X vssd1 vssd1 vccd1 vccd1 _09168_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08119_ _09541_/C _07974_/B _08118_/X vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__o21ai_1
X_09099_ _15558_/Q _09220_/B _09099_/C vssd1 vssd1 vccd1 vccd1 _09101_/C sky130_fd_sc_hd__nand3_1
X_11130_ _11123_/C _11124_/C _11126_/Y _11128_/X vssd1 vssd1 vccd1 vccd1 _11131_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11061_ _15919_/Q _11118_/B _11070_/C vssd1 vssd1 vccd1 vccd1 _11066_/A sky130_fd_sc_hd__and3_1
X_10012_ _10716_/A vssd1 vssd1 vccd1 vccd1 _10012_/X sky130_fd_sc_hd__buf_2
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14820_ _14820_/A vssd1 vssd1 vccd1 vccd1 _16456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14751_ _14747_/Y _14748_/X _14750_/Y _14745_/C vssd1 vssd1 vccd1 vccd1 _14753_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11963_ _11963_/A vssd1 vssd1 vccd1 vccd1 _12084_/A sky130_fd_sc_hd__buf_2
XFILLER_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13702_ _13699_/Y _13711_/A _13701_/Y _13696_/C vssd1 vssd1 vccd1 vccd1 _13704_/B
+ sky130_fd_sc_hd__o211a_1
X_10914_ _15897_/Q _11026_/B _10914_/C vssd1 vssd1 vccd1 vccd1 _10914_/Y sky130_fd_sc_hd__nand3_1
XFILLER_72_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11894_ _11892_/Y _11888_/C _11890_/Y _11899_/A vssd1 vssd1 vccd1 vccd1 _11899_/B
+ sky130_fd_sc_hd__a211oi_1
X_14682_ _16436_/Q _14689_/C _14567_/X vssd1 vssd1 vccd1 vccd1 _14685_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16421_ _16595_/CLK _16421_/D vssd1 vssd1 vccd1 vccd1 _16421_/Q sky130_fd_sc_hd__dfxtp_1
X_10845_ _10841_/Y _10844_/X _10838_/C _10839_/C vssd1 vssd1 vccd1 vccd1 _10847_/B
+ sky130_fd_sc_hd__o211ai_1
X_13633_ _13630_/Y _13631_/X _13632_/Y _13628_/C vssd1 vssd1 vccd1 vccd1 _13635_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16352_ _16389_/CLK _16352_/D vssd1 vssd1 vccd1 vccd1 _16352_/Q sky130_fd_sc_hd__dfxtp_1
X_13564_ _16273_/Q _13573_/C _13450_/X vssd1 vssd1 vccd1 vccd1 _13564_/Y sky130_fd_sc_hd__a21oi_1
X_10776_ _10777_/B _10777_/C _10777_/A vssd1 vssd1 vccd1 vccd1 _10778_/B sky130_fd_sc_hd__a21o_1
X_15303_ _15303_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15304_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12515_ _16125_/Q _12516_/C _12292_/X vssd1 vssd1 vccd1 vccd1 _12517_/A sky130_fd_sc_hd__a21oi_1
X_13495_ _14060_/A vssd1 vssd1 vccd1 vccd1 _13495_/X sky130_fd_sc_hd__clkbuf_2
X_16283_ _16346_/CLK _16283_/D vssd1 vssd1 vccd1 vccd1 _16283_/Q sky130_fd_sc_hd__dfxtp_1
X_15234_ _16526_/Q _15241_/C _10956_/A vssd1 vssd1 vccd1 vccd1 _15237_/B sky130_fd_sc_hd__a21o_1
X_12446_ _12453_/A _12446_/B _12446_/C vssd1 vssd1 vccd1 vccd1 _12447_/A sky130_fd_sc_hd__and3_1
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15165_ _15271_/A _15169_/C vssd1 vssd1 vccd1 vccd1 _15165_/X sky130_fd_sc_hd__or2_1
X_12377_ _12398_/A _12377_/B _12377_/C vssd1 vssd1 vccd1 vccd1 _12378_/A sky130_fd_sc_hd__and3_1
XFILLER_126_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11328_ _15957_/Q _11381_/B _11328_/C vssd1 vssd1 vccd1 vccd1 _11336_/B sky130_fd_sc_hd__and3_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ _14148_/C vssd1 vssd1 vccd1 vccd1 _14154_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15096_ _16502_/Q _15254_/B _15103_/C vssd1 vssd1 vccd1 vccd1 _15096_/X sky130_fd_sc_hd__and3_1
XFILLER_140_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11259_ _15947_/Q _11367_/B _11268_/C vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__and3_1
X_14047_ _14047_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14053_/C sky130_fd_sc_hd__nor2_1
XFILLER_140_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15998_ _16005_/CLK _15998_/D vssd1 vssd1 vccd1 vccd1 _15998_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ _14949_/A _14949_/B vssd1 vssd1 vccd1 vccd1 _14950_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08470_ _08403_/A _08403_/B _08469_/Y vssd1 vssd1 vccd1 vccd1 _08512_/B sky130_fd_sc_hd__a21oi_4
XFILLER_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16619_ input11/X _16619_/D vssd1 vssd1 vccd1 vccd1 _16619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09022_ _15541_/Q _09145_/B _09028_/C vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__and3_1
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09924_ _09921_/A _09920_/Y _09921_/B vssd1 vssd1 vccd1 vccd1 _09924_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_120_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _10276_/A vssd1 vssd1 vccd1 vccd1 _09855_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _15495_/Q _08807_/C _08805_/X vssd1 vssd1 vccd1 vccd1 _08809_/B sky130_fd_sc_hd__a21o_1
X_09786_ _09780_/Y _09781_/X _09783_/B vssd1 vssd1 vccd1 vccd1 _09787_/B sky130_fd_sc_hd__o21a_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08737_ _08735_/A _08735_/B _08736_/X vssd1 vssd1 vccd1 vccd1 _15475_/D sky130_fd_sc_hd__a21oi_1
XFILLER_39_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _16551_/Q _16550_/Q _16549_/Q _08667_/X vssd1 vssd1 vccd1 vccd1 _15462_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ input2/X vssd1 vssd1 vccd1 vccd1 _12886_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_121_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10630_ _15852_/Q _10726_/B _10630_/C vssd1 vssd1 vccd1 vccd1 _10635_/A sky130_fd_sc_hd__and3_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10561_ _10558_/Y _10567_/A _10560_/Y _10556_/C vssd1 vssd1 vccd1 vccd1 _10563_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12300_ _12466_/A _12304_/C vssd1 vssd1 vccd1 vccd1 _12300_/X sky130_fd_sc_hd__or2_1
XFILLER_10_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13280_ _13302_/A _13280_/B _13280_/C vssd1 vssd1 vccd1 vccd1 _13281_/A sky130_fd_sc_hd__and3_1
X_10492_ _10492_/A vssd1 vssd1 vccd1 vccd1 _10492_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ _16085_/Q _12232_/C _12007_/X vssd1 vssd1 vccd1 vccd1 _12233_/A sky130_fd_sc_hd__a21oi_1
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12162_ _12160_/Y _12155_/C _12158_/Y _12159_/X vssd1 vssd1 vccd1 vccd1 _12163_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11113_ _11113_/A vssd1 vssd1 vccd1 vccd1 _11128_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12093_ _16065_/Q _12204_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__and3_1
XFILLER_77_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11044_ _15917_/Q _11045_/C _10874_/X vssd1 vssd1 vccd1 vccd1 _11046_/A sky130_fd_sc_hd__a21oi_1
X_15921_ _16005_/CLK _15921_/D vssd1 vssd1 vccd1 vccd1 _15921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15852_ _16595_/CLK _15852_/D vssd1 vssd1 vccd1 vccd1 _15852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14803_ _14819_/A _14803_/B _14803_/C vssd1 vssd1 vccd1 vccd1 _14804_/A sky130_fd_sc_hd__and3_1
X_15783_ _15812_/CLK _15783_/D vssd1 vssd1 vccd1 vccd1 _15783_/Q sky130_fd_sc_hd__dfxtp_1
X_12995_ _16192_/Q _13164_/B _13001_/C vssd1 vssd1 vccd1 vccd1 _12997_/C sky130_fd_sc_hd__nand3_1
XFILLER_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14734_ _14768_/A _14734_/B _14738_/A vssd1 vssd1 vccd1 vccd1 _16443_/D sky130_fd_sc_hd__nor3_1
X_11946_ _11942_/Y _11952_/A _11945_/Y _11940_/C vssd1 vssd1 vccd1 vccd1 _11948_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14665_ _14665_/A _14665_/B vssd1 vssd1 vccd1 vccd1 _14671_/C sky130_fd_sc_hd__nor2_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ _16034_/Q _11928_/B _11878_/C vssd1 vssd1 vccd1 vccd1 _11877_/X sky130_fd_sc_hd__and3_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16404_ _16607_/CLK _16404_/D vssd1 vssd1 vccd1 vccd1 _16404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13616_ _16281_/Q _13625_/C _13450_/X vssd1 vssd1 vccd1 vccd1 _13616_/Y sky130_fd_sc_hd__a21oi_1
X_10828_ _16557_/Q vssd1 vssd1 vccd1 vccd1 _10844_/C sky130_fd_sc_hd__inv_2
X_14596_ _16422_/Q _14603_/C _14537_/X vssd1 vssd1 vccd1 vccd1 _14596_/Y sky130_fd_sc_hd__a21oi_1
X_16335_ _16346_/CLK _16335_/D vssd1 vssd1 vccd1 vccd1 _16335_/Q sky130_fd_sc_hd__dfxtp_1
X_13547_ _13548_/B _13548_/C _13546_/X vssd1 vssd1 vccd1 vccd1 _13549_/B sky130_fd_sc_hd__o21ai_1
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10759_ _10759_/A _10759_/B vssd1 vssd1 vccd1 vccd1 _10759_/X sky130_fd_sc_hd__or2_1
X_16266_ _16533_/Q _16266_/D vssd1 vssd1 vccd1 vccd1 _16266_/Q sky130_fd_sc_hd__dfxtp_1
X_13478_ _16261_/Q _13479_/C _13421_/X vssd1 vssd1 vccd1 vccd1 _13480_/A sky130_fd_sc_hd__a21oi_1
XFILLER_145_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15217_ _15217_/A _15217_/B vssd1 vssd1 vccd1 vccd1 _15218_/B sky130_fd_sc_hd__nor2_1
X_12429_ _16112_/Q _12600_/B _12435_/C vssd1 vssd1 vccd1 vccd1 _12431_/C sky130_fd_sc_hd__nand3_1
X_16197_ _16555_/Q _16197_/D vssd1 vssd1 vccd1 vccd1 _16197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15148_ _16511_/Q _15254_/B _15155_/C vssd1 vssd1 vccd1 vccd1 _15148_/X sky130_fd_sc_hd__and3_1
XFILLER_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07970_ _10675_/C _07970_/B vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__xnor2_1
XFILLER_141_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15079_ _15079_/A _15079_/B _15079_/C vssd1 vssd1 vccd1 vccd1 _15080_/C sky130_fd_sc_hd__nand3_1
XFILLER_101_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09640_ _15667_/Q _09648_/C _09463_/X vssd1 vssd1 vccd1 vccd1 _09643_/A sky130_fd_sc_hd__a21oi_1
XFILLER_68_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ _09529_/X _09568_/B _09570_/Y vssd1 vssd1 vccd1 vccd1 _15649_/D sky130_fd_sc_hd__o21a_1
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08522_ _15451_/Q _08561_/B _15307_/C vssd1 vssd1 vccd1 vccd1 _08564_/A sky130_fd_sc_hd__and3_1
XFILLER_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08453_ _08453_/A _08505_/A vssd1 vssd1 vccd1 vccd1 _08496_/A sky130_fd_sc_hd__xnor2_4
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08384_ _08384_/A _08455_/A vssd1 vssd1 vccd1 vccd1 _08395_/A sky130_fd_sc_hd__xnor2_4
XFILLER_109_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09005_ _09005_/A _09005_/B vssd1 vssd1 vccd1 vccd1 _15532_/D sky130_fd_sc_hd__nor2_1
XFILLER_132_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09907_ _15719_/Q _09914_/C _08589_/A vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09838_ _15702_/Q _10308_/C _09845_/C vssd1 vssd1 vccd1 vccd1 _09838_/Y sky130_fd_sc_hd__nand3_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16682__87 vssd1 vssd1 vccd1 vccd1 _16682__87/HI _16758_/A sky130_fd_sc_hd__conb_1
XFILLER_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09769_ _15693_/Q _09770_/C _09590_/X vssd1 vssd1 vccd1 vccd1 _09769_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _11821_/C vssd1 vssd1 vccd1 vccd1 _11836_/C sky130_fd_sc_hd__clkbuf_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12778_/Y _12773_/C _12775_/Y _12776_/X vssd1 vssd1 vccd1 vccd1 _12781_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _11731_/A _11731_/B vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__nor2_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14484_/A _14450_/B _14454_/A vssd1 vssd1 vccd1 vccd1 _16398_/D sky130_fd_sc_hd__nor3_1
XFILLER_30_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11662_ _16004_/Q _11891_/B _11662_/C vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__and3_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13401_ _16249_/Q _13573_/B _13401_/C vssd1 vssd1 vccd1 vccd1 _13401_/Y sky130_fd_sc_hd__nand3_1
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10613_ _10613_/A _10613_/B vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__or2_1
X_11593_ _15994_/Q _11644_/B _11594_/C vssd1 vssd1 vccd1 vccd1 _11593_/X sky130_fd_sc_hd__and3_1
X_14381_ _14381_/A _14389_/B vssd1 vssd1 vccd1 vccd1 _14383_/A sky130_fd_sc_hd__or2_1
X_16120_ _16554_/Q _16120_/D vssd1 vssd1 vccd1 vccd1 _16120_/Q sky130_fd_sc_hd__dfxtp_1
X_13332_ _13332_/A _13332_/B _13332_/C vssd1 vssd1 vccd1 vccd1 _13333_/C sky130_fd_sc_hd__nand3_1
X_10544_ _15836_/Q _10546_/C _10492_/X vssd1 vssd1 vccd1 vccd1 _10544_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16051_ _16118_/CLK _16051_/D vssd1 vssd1 vccd1 vccd1 _16051_/Q sky130_fd_sc_hd__dfxtp_1
X_10475_ _10276_/X _10471_/B _10474_/Y vssd1 vssd1 vccd1 vccd1 _15821_/D sky130_fd_sc_hd__o21a_1
X_13263_ _13317_/A vssd1 vssd1 vccd1 vccd1 _13302_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15002_ _15002_/A _15009_/B vssd1 vssd1 vccd1 vccd1 _15004_/A sky130_fd_sc_hd__or2_1
X_12214_ _12212_/Y _12207_/C _12209_/Y _12210_/X vssd1 vssd1 vccd1 vccd1 _12215_/C
+ sky130_fd_sc_hd__a211o_1
X_13194_ _16219_/Q _13194_/B _13199_/C vssd1 vssd1 vccd1 vccd1 _13194_/Y sky130_fd_sc_hd__nand3_1
X_12145_ _16072_/Q _12152_/C _12029_/X vssd1 vssd1 vccd1 vccd1 _12148_/B sky130_fd_sc_hd__a21o_1
XFILLER_150_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12076_ _12076_/A vssd1 vssd1 vccd1 vccd1 _16061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ _11024_/Y _11025_/X _11026_/Y _11021_/C vssd1 vssd1 vccd1 vccd1 _11029_/B
+ sky130_fd_sc_hd__o211ai_1
X_15904_ _16553_/Q _15904_/D vssd1 vssd1 vccd1 vccd1 _15904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15835_ _16570_/CLK _15835_/D vssd1 vssd1 vccd1 vccd1 _15835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15766_ _15812_/CLK _15766_/D vssd1 vssd1 vccd1 vccd1 _15766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _12978_/A _12978_/B vssd1 vssd1 vccd1 vccd1 _12984_/C sky130_fd_sc_hd__nor2_1
XFILLER_17_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14717_ _14717_/A _14724_/B vssd1 vssd1 vccd1 vccd1 _14719_/A sky130_fd_sc_hd__or2_1
X_11929_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12160_/B sky130_fd_sc_hd__clkbuf_2
X_15697_ _15791_/CLK _15697_/D vssd1 vssd1 vccd1 vccd1 _15697_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14648_ _16429_/Q _14875_/B _14655_/C vssd1 vssd1 vccd1 vccd1 _14648_/Y sky130_fd_sc_hd__nand3_1
XFILLER_14_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_17 _11384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _09125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14579_ _14594_/A _14579_/B _14579_/C vssd1 vssd1 vccd1 vccd1 _14580_/A sky130_fd_sc_hd__and3_1
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16318_ _16346_/CLK _16318_/D vssd1 vssd1 vccd1 vccd1 _16318_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16249_ _16261_/CLK _16249_/D vssd1 vssd1 vccd1 vccd1 _16249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07953_ _16576_/Q vssd1 vssd1 vccd1 vccd1 _11908_/A sky130_fd_sc_hd__inv_2
X_07884_ _16618_/Q vssd1 vssd1 vccd1 vccd1 _14279_/A sky130_fd_sc_hd__inv_2
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09623_ _09636_/C vssd1 vssd1 vccd1 vccd1 _09648_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09554_ _15649_/Q _09561_/C _09463_/X vssd1 vssd1 vccd1 vccd1 _09557_/A sky130_fd_sc_hd__a21oi_1
XFILLER_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08505_ _08505_/A _08453_/A vssd1 vssd1 vccd1 vccd1 _08509_/B sky130_fd_sc_hd__or2b_1
XFILLER_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09485_ _09394_/X _09481_/B _09351_/X vssd1 vssd1 vccd1 vccd1 _09489_/A sky130_fd_sc_hd__a21oi_1
XFILLER_63_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08436_ _08343_/A _08343_/B _08435_/Y vssd1 vssd1 vccd1 vccd1 _08446_/A sky130_fd_sc_hd__a21o_2
XFILLER_11_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08367_ _08367_/A _08437_/A vssd1 vssd1 vccd1 vccd1 _08403_/A sky130_fd_sc_hd__xnor2_4
X_08298_ _08298_/A _08299_/A vssd1 vssd1 vccd1 vccd1 _08300_/A sky130_fd_sc_hd__or2b_1
XFILLER_137_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10260_ _15784_/Q _10267_/C _10204_/X vssd1 vssd1 vccd1 vccd1 _10260_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10191_ _10189_/Y _10190_/X _10186_/C _10187_/C vssd1 vssd1 vccd1 vccd1 _10193_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_87_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13950_ _16328_/Q _13958_/C _13729_/X vssd1 vssd1 vccd1 vccd1 _13953_/B sky130_fd_sc_hd__a21o_1
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12901_ _12901_/A vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__buf_2
X_13881_ _13881_/A vssd1 vssd1 vccd1 vccd1 _13918_/A sky130_fd_sc_hd__clkbuf_2
X_15620_ _15812_/CLK _15620_/D vssd1 vssd1 vccd1 vccd1 _15620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12832_ _12832_/A vssd1 vssd1 vccd1 vccd1 _16168_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15551_ _16551_/CLK _15551_/D vssd1 vssd1 vccd1 vccd1 _15551_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _16160_/Q _12770_/C _12598_/X vssd1 vssd1 vccd1 vccd1 _12766_/B sky130_fd_sc_hd__a21o_1
XFILLER_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14516_/C vssd1 vssd1 vccd1 vccd1 _14524_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _16010_/Q _11773_/B _11721_/C vssd1 vssd1 vccd1 vccd1 _11714_/Y sky130_fd_sc_hd__nand3_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _16570_/CLK _15482_/D vssd1 vssd1 vccd1 vccd1 _15482_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12694_/A _12694_/B vssd1 vssd1 vccd1 vccd1 _12695_/B sky130_fd_sc_hd__nor2_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _16397_/Q _14486_/B _14433_/C vssd1 vssd1 vccd1 vccd1 _14441_/B sky130_fd_sc_hd__and3_1
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11645_ _12886_/A vssd1 vssd1 vccd1 vccd1 _15241_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14364_ _16387_/Q _14472_/B _14373_/C vssd1 vssd1 vccd1 vccd1 _14364_/X sky130_fd_sc_hd__and3_1
X_11576_ _15991_/Q _11613_/C _11517_/X vssd1 vssd1 vccd1 vccd1 _11578_/B sky130_fd_sc_hd__a21oi_1
XFILLER_6_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16103_ _16118_/CLK _16103_/D vssd1 vssd1 vccd1 vccd1 _16103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13315_ _13315_/A _13319_/C vssd1 vssd1 vccd1 vccd1 _13315_/X sky130_fd_sc_hd__or2_1
X_10527_ _10418_/X _10524_/B _10473_/X vssd1 vssd1 vccd1 vccd1 _10527_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14295_ _16377_/Q _14303_/C _14294_/X vssd1 vssd1 vccd1 vccd1 _14295_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_143_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16034_ _16118_/CLK _16034_/D vssd1 vssd1 vccd1 vccd1 _16034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10458_ _15819_/Q _10458_/B _10463_/C vssd1 vssd1 vccd1 vccd1 _10458_/Y sky130_fd_sc_hd__nand3_1
X_13246_ _13246_/A _13246_/B _13246_/C vssd1 vssd1 vccd1 vccd1 _13247_/A sky130_fd_sc_hd__and3_1
XFILLER_124_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ _10387_/Y _10388_/X _10384_/C _10385_/C vssd1 vssd1 vccd1 vccd1 _10391_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_123_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13177_ _16218_/Q _13342_/B _13178_/C vssd1 vssd1 vccd1 vccd1 _13177_/X sky130_fd_sc_hd__and3_1
XFILLER_111_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12128_ _12128_/A _12128_/B vssd1 vssd1 vccd1 vccd1 _12135_/C sky130_fd_sc_hd__nor2_1
XFILLER_97_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12059_ _16060_/Q _12173_/B _12059_/C vssd1 vssd1 vccd1 vccd1 _12067_/A sky130_fd_sc_hd__and3_1
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15818_ _16570_/CLK _15818_/D vssd1 vssd1 vccd1 vccd1 _15818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15749_ _15812_/CLK _15749_/D vssd1 vssd1 vccd1 vccd1 _15749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09270_ _09374_/A _09270_/B _09276_/B vssd1 vssd1 vccd1 vccd1 _15591_/D sky130_fd_sc_hd__nor3_1
XFILLER_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08221_ _08373_/B _08454_/B vssd1 vssd1 vccd1 vccd1 _08368_/A sky130_fd_sc_hd__xor2_4
XFILLER_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08152_ _13322_/A _07912_/B _08151_/X vssd1 vssd1 vccd1 vccd1 _08160_/A sky130_fd_sc_hd__o21ai_1
X_08083_ _08254_/A _08083_/B vssd1 vssd1 vccd1 vccd1 _08088_/A sky130_fd_sc_hd__xnor2_4
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08985_ _15532_/Q _09145_/B _08991_/C vssd1 vssd1 vccd1 vccd1 _08993_/A sky130_fd_sc_hd__and3_1
XFILLER_102_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07936_ _16534_/Q _16532_/Q vssd1 vssd1 vccd1 vccd1 _08265_/A sky130_fd_sc_hd__nand2_2
X_07867_ _16594_/Q vssd1 vssd1 vccd1 vccd1 _12928_/A sky130_fd_sc_hd__inv_2
X_16652__57 vssd1 vssd1 vccd1 vccd1 _16652__57/HI _16728_/A sky130_fd_sc_hd__conb_1
XFILLER_113_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _09603_/X _09606_/B vssd1 vssd1 vccd1 vccd1 _09606_/X sky130_fd_sc_hd__and2b_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07798_ _07799_/A vssd1 vssd1 vccd1 vccd1 _07798_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09537_ _15632_/Q _15631_/Q _15630_/Q _09536_/X vssd1 vssd1 vccd1 vccd1 _15642_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _09468_/A _09468_/B vssd1 vssd1 vccd1 vccd1 _09468_/X sky130_fd_sc_hd__or2_1
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08419_ _08419_/A _08419_/B vssd1 vssd1 vccd1 vccd1 _08419_/X sky130_fd_sc_hd__and2_1
X_09399_ _15605_/Q _15604_/Q _15603_/Q _09314_/X vssd1 vssd1 vccd1 vccd1 _15615_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11430_ _11428_/Y _11423_/C _11425_/Y _11427_/X vssd1 vssd1 vccd1 vccd1 _11431_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _15961_/Q _11594_/B _11361_/C vssd1 vssd1 vccd1 vccd1 _11361_/Y sky130_fd_sc_hd__nand3_1
XFILLER_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10312_ _15794_/Q _10313_/B _10104_/X vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__a21oi_1
X_13100_ _13135_/C vssd1 vssd1 vccd1 vccd1 _13143_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11292_ _15951_/Q _11402_/B _11301_/C vssd1 vssd1 vccd1 vccd1 _11297_/A sky130_fd_sc_hd__and3_1
X_14080_ _14077_/Y _14078_/X _14079_/Y _14075_/C vssd1 vssd1 vccd1 vccd1 _14082_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10243_ _10492_/A vssd1 vssd1 vccd1 vccd1 _10243_/X sky130_fd_sc_hd__buf_2
X_13031_ _13031_/A _13031_/B vssd1 vssd1 vccd1 vccd1 _13036_/C sky130_fd_sc_hd__nor2_1
XFILLER_106_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10174_ _10206_/C vssd1 vssd1 vccd1 vccd1 _10214_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_78_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14982_ _16482_/Q _14982_/B _14982_/C vssd1 vssd1 vccd1 vccd1 _14982_/Y sky130_fd_sc_hd__nand3_1
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16721_ _16721_/A _07826_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
XFILLER_87_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13933_ _13933_/A _13933_/B vssd1 vssd1 vccd1 vccd1 _13939_/C sky130_fd_sc_hd__nor2_1
XFILLER_35_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13864_ _13861_/Y _13862_/X _13863_/Y _13859_/C vssd1 vssd1 vccd1 vccd1 _13866_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_28_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15603_ _16551_/CLK _15603_/D vssd1 vssd1 vccd1 vccd1 _15603_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ _12836_/C vssd1 vssd1 vccd1 vccd1 _12852_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16583_ _16595_/CLK _16583_/D vssd1 vssd1 vccd1 vccd1 _16583_/Q sky130_fd_sc_hd__dfxtp_1
X_13795_ _13789_/C _13790_/C _13792_/Y _13793_/X vssd1 vssd1 vccd1 vccd1 _13796_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15534_ _16551_/CLK _15534_/D vssd1 vssd1 vccd1 vccd1 _15534_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _12746_/A _12753_/B vssd1 vssd1 vccd1 vccd1 _12748_/A sky130_fd_sc_hd__or2_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15465_ _16570_/CLK _15465_/D vssd1 vssd1 vccd1 vccd1 _15465_/Q sky130_fd_sc_hd__dfxtp_2
X_12677_ _13242_/A vssd1 vssd1 vccd1 vccd1 _12904_/B sky130_fd_sc_hd__buf_2
XFILLER_147_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14416_ _14414_/Y _14409_/C _14412_/Y _14413_/X vssd1 vssd1 vccd1 vccd1 _14417_/C
+ sky130_fd_sc_hd__a211o_1
X_11628_ _15999_/Q _11668_/C _11517_/X vssd1 vssd1 vccd1 vccd1 _11630_/B sky130_fd_sc_hd__a21oi_1
X_15396_ _16069_/Q _16068_/Q _16067_/Q _15391_/X vssd1 vssd1 vccd1 vccd1 _16579_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14347_ _14347_/A _14347_/B _14347_/C vssd1 vssd1 vccd1 vccd1 _14348_/C sky130_fd_sc_hd__nand3_1
XFILLER_129_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11559_ _15989_/Q _11560_/C _11441_/X vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__a21oi_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ _14278_/A vssd1 vssd1 vccd1 vccd1 _16373_/D sky130_fd_sc_hd__clkbuf_1
X_16017_ _16554_/Q _16017_/D vssd1 vssd1 vccd1 vccd1 _16017_/Q sky130_fd_sc_hd__dfxtp_1
X_13229_ _13227_/Y _13228_/X _13224_/C _13225_/C vssd1 vssd1 vccd1 vccd1 _13231_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _08770_/A vssd1 vssd1 vccd1 vccd1 _15482_/D sky130_fd_sc_hd__clkbuf_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09322_ _15602_/Q _09329_/C _09992_/B vssd1 vssd1 vccd1 vccd1 _09325_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09253_ _15592_/Q _09286_/C _09252_/X vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08204_ _08204_/A _08204_/B _08204_/C vssd1 vssd1 vccd1 vccd1 _08205_/B sky130_fd_sc_hd__and3_1
X_09184_ _10294_/C vssd1 vssd1 vccd1 vccd1 _15341_/B sky130_fd_sc_hd__clkbuf_4
X_08135_ _08135_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _08325_/A sky130_fd_sc_hd__xnor2_4
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08066_ _14785_/A _08066_/B vssd1 vssd1 vccd1 vccd1 _08245_/B sky130_fd_sc_hd__xnor2_2
XFILLER_135_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08968_ _15515_/Q _15514_/Q _15513_/Q _08887_/X vssd1 vssd1 vccd1 vccd1 _15525_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07919_ _16606_/Q vssd1 vssd1 vccd1 vccd1 _13603_/A sky130_fd_sc_hd__clkinv_2
XFILLER_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08899_ _08940_/A _08899_/B _08899_/C vssd1 vssd1 vccd1 vccd1 _08900_/A sky130_fd_sc_hd__and3_1
X_10930_ _10927_/Y _10936_/A _10929_/Y _10925_/C vssd1 vssd1 vccd1 vccd1 _10932_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861_ _15890_/Q _10922_/B _10868_/C vssd1 vssd1 vccd1 vccd1 _10861_/Y sky130_fd_sc_hd__nand3_1
XFILLER_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12600_ _16136_/Q _12600_/B _12607_/C vssd1 vssd1 vccd1 vccd1 _12602_/C sky130_fd_sc_hd__nand3_1
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _16274_/Q _13753_/B _13586_/C vssd1 vssd1 vccd1 vccd1 _13580_/Y sky130_fd_sc_hd__nand3_1
XFILLER_25_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10792_ _10788_/Y _10789_/X _10791_/Y _10785_/C vssd1 vssd1 vccd1 vccd1 _10794_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12545_/C vssd1 vssd1 vccd1 vccd1 _12554_/C sky130_fd_sc_hd__clkbuf_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15250_ _15248_/Y _15244_/C _15246_/Y _15247_/X vssd1 vssd1 vccd1 vccd1 _15251_/C
+ sky130_fd_sc_hd__a211o_1
X_12462_ _16117_/Q _12516_/B _12462_/C vssd1 vssd1 vccd1 vccd1 _12470_/B sky130_fd_sc_hd__and3_1
X_14201_ _16364_/Q _14427_/B _14201_/C vssd1 vssd1 vccd1 vccd1 _14209_/A sky130_fd_sc_hd__and3_1
XFILLER_138_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11413_ _11410_/Y _11412_/X _11407_/C _11408_/C vssd1 vssd1 vccd1 vccd1 _11415_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_149_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15181_ _16517_/Q _15188_/C _10956_/A vssd1 vssd1 vccd1 vccd1 _15184_/B sky130_fd_sc_hd__a21o_1
X_12393_ _16107_/Q _12501_/B _12402_/C vssd1 vssd1 vccd1 vccd1 _12393_/X sky130_fd_sc_hd__and3_1
XFILLER_125_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14132_ _14411_/A vssd1 vssd1 vccd1 vccd1 _14132_/X sky130_fd_sc_hd__clkbuf_2
X_11344_ _15959_/Q _11402_/B _11353_/C vssd1 vssd1 vccd1 vccd1 _11349_/A sky130_fd_sc_hd__and3_1
XFILLER_4_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14063_ _14063_/A _14063_/B _14068_/A vssd1 vssd1 vccd1 vccd1 _16342_/D sky130_fd_sc_hd__nor3_1
X_11275_ _15949_/Q _11381_/B _11275_/C vssd1 vssd1 vccd1 vccd1 _11284_/B sky130_fd_sc_hd__and3_1
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13014_ _16195_/Q _13022_/C _12901_/X vssd1 vssd1 vccd1 vccd1 _13014_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10226_ _09855_/X _10222_/B _10225_/Y vssd1 vssd1 vccd1 vccd1 _15776_/D sky130_fd_sc_hd__o21a_1
XFILLER_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10157_ _15767_/Q _10158_/C _10104_/X vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__a21oi_1
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10088_ _10081_/C _10082_/C _10085_/Y _10086_/X vssd1 vssd1 vccd1 vccd1 _10089_/C
+ sky130_fd_sc_hd__a211o_1
X_14965_ _16480_/Q _15074_/B _14974_/C vssd1 vssd1 vccd1 vccd1 _14970_/A sky130_fd_sc_hd__and3_1
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16704_ _16704_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13916_ _13913_/Y _13914_/X _13915_/Y _13911_/C vssd1 vssd1 vccd1 vccd1 _13918_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14896_ _15117_/A _14896_/B _14896_/C vssd1 vssd1 vccd1 vccd1 _14897_/C sky130_fd_sc_hd__or3_1
XFILLER_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13847_ _16313_/Q _13856_/C _13736_/X vssd1 vssd1 vccd1 vccd1 _13847_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16566_ _16570_/CLK _16566_/D vssd1 vssd1 vccd1 vccd1 _16566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13778_ _13793_/C vssd1 vssd1 vccd1 vccd1 _13800_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15517_ _15791_/CLK _15517_/D vssd1 vssd1 vccd1 vccd1 _15517_/Q sky130_fd_sc_hd__dfxtp_2
X_12729_ _12736_/A _12729_/B _12729_/C vssd1 vssd1 vccd1 vccd1 _12730_/A sky130_fd_sc_hd__and3_1
X_16497_ _16607_/CLK _16497_/D vssd1 vssd1 vccd1 vccd1 _16497_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15448_ _16570_/CLK _15448_/D vssd1 vssd1 vccd1 vccd1 _15448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15379_ _15957_/Q _15956_/Q _15955_/Q _15378_/X vssd1 vssd1 vccd1 vccd1 _16565_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_128_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09940_ _15741_/Q vssd1 vssd1 vccd1 vccd1 _09945_/C sky130_fd_sc_hd__inv_2
XFILLER_143_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _09871_/A vssd1 vssd1 vccd1 vccd1 _15707_/D sky130_fd_sc_hd__clkbuf_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _15497_/Q _08991_/B _08822_/C vssd1 vssd1 vccd1 vccd1 _08823_/B sky130_fd_sc_hd__and3_1
XFILLER_98_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _08706_/X _08745_/A _08708_/X vssd1 vssd1 vccd1 vccd1 _08754_/B sky130_fd_sc_hd__o21ai_1
XFILLER_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _15469_/Q _10743_/B _08689_/C vssd1 vssd1 vccd1 vccd1 _08691_/A sky130_fd_sc_hd__and3_1
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16622__27 vssd1 vssd1 vccd1 vccd1 _16622__27/HI _16688_/A sky130_fd_sc_hd__conb_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ _09301_/X _09296_/B _09304_/X vssd1 vssd1 vccd1 vccd1 _09305_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09236_ _09234_/A _09234_/B _09235_/X vssd1 vssd1 vccd1 vccd1 _15583_/D sky130_fd_sc_hd__a21oi_1
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09167_ _09167_/A _09167_/B vssd1 vssd1 vccd1 vccd1 _15568_/D sky130_fd_sc_hd__nor2_1
X_08118_ _09625_/C _08118_/B vssd1 vssd1 vccd1 vccd1 _08118_/X sky130_fd_sc_hd__or2_1
XFILLER_134_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _15558_/Q _09099_/C _09014_/X vssd1 vssd1 vccd1 vccd1 _09101_/B sky130_fd_sc_hd__a21o_1
XFILLER_79_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08049_ _14559_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08229_/B sky130_fd_sc_hd__xnor2_4
XFILLER_122_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11060_ _15919_/Q _11099_/C _10951_/X vssd1 vssd1 vccd1 vccd1 _11062_/B sky130_fd_sc_hd__a21oi_1
X_10011_ _10009_/X _10011_/B vssd1 vssd1 vccd1 vccd1 _10011_/X sky130_fd_sc_hd__and2b_1
XFILLER_89_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14750_ _16446_/Q _14982_/B _14750_/C vssd1 vssd1 vccd1 vccd1 _14750_/Y sky130_fd_sc_hd__nand3_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11962_ _11962_/A vssd1 vssd1 vccd1 vccd1 _16045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13701_ _16291_/Q _13760_/B _13709_/C vssd1 vssd1 vccd1 vccd1 _13701_/Y sky130_fd_sc_hd__nand3_1
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10913_ _15898_/Q _11076_/B _10914_/C vssd1 vssd1 vccd1 vccd1 _10913_/X sky130_fd_sc_hd__and3_1
X_14681_ _14768_/A _14681_/B _14685_/A vssd1 vssd1 vccd1 vccd1 _16434_/D sky130_fd_sc_hd__nor3_1
X_11893_ _11890_/Y _11899_/A _11892_/Y _11888_/C vssd1 vssd1 vccd1 vccd1 _11895_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16420_ _16595_/CLK _16420_/D vssd1 vssd1 vccd1 vccd1 _16420_/Q sky130_fd_sc_hd__dfxtp_1
X_13632_ _16282_/Q _13753_/B _13639_/C vssd1 vssd1 vccd1 vccd1 _13632_/Y sky130_fd_sc_hd__nand3_1
XFILLER_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ _15889_/Q _11070_/B _10844_/C vssd1 vssd1 vccd1 vccd1 _10844_/X sky130_fd_sc_hd__and3_1
X_16351_ _16389_/CLK _16351_/D vssd1 vssd1 vccd1 vccd1 _16351_/Q sky130_fd_sc_hd__dfxtp_1
X_13563_ _13563_/A vssd1 vssd1 vccd1 vccd1 _16271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10775_ _15879_/Q _10900_/B _10782_/C vssd1 vssd1 vccd1 vccd1 _10777_/C sky130_fd_sc_hd__nand3_1
X_15302_ _15292_/A _15294_/X _15292_/B vssd1 vssd1 vccd1 vccd1 _15303_/B sky130_fd_sc_hd__a21bo_1
X_12514_ _12514_/A _12514_/B _12518_/B vssd1 vssd1 vccd1 vccd1 _16123_/D sky130_fd_sc_hd__nor3_1
X_16282_ _16533_/Q _16282_/D vssd1 vssd1 vccd1 vccd1 _16282_/Q sky130_fd_sc_hd__dfxtp_1
X_13494_ _13531_/C vssd1 vssd1 vccd1 vccd1 _13538_/C sky130_fd_sc_hd__clkbuf_2
X_15233_ _15333_/A _15233_/B _15237_/A vssd1 vssd1 vccd1 vccd1 _16524_/D sky130_fd_sc_hd__nor3_1
X_12445_ _12443_/Y _12438_/C _12441_/Y _12442_/X vssd1 vssd1 vccd1 vccd1 _12446_/C
+ sky130_fd_sc_hd__a211o_1
X_15164_ _15164_/A _15164_/B vssd1 vssd1 vccd1 vccd1 _15169_/C sky130_fd_sc_hd__nor2_1
X_12376_ _12376_/A _12376_/B _12376_/C vssd1 vssd1 vccd1 vccd1 _12377_/C sky130_fd_sc_hd__nand3_1
XFILLER_125_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14115_ _14135_/C vssd1 vssd1 vccd1 vccd1 _14148_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11327_ _15957_/Q _11328_/C _11158_/X vssd1 vssd1 vccd1 vccd1 _11329_/A sky130_fd_sc_hd__a21oi_1
XFILLER_114_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15095_ _16502_/Q _15103_/C _14872_/X vssd1 vssd1 vccd1 vccd1 _15095_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14046_ _14046_/A _14046_/B vssd1 vssd1 vccd1 vccd1 _14047_/B sky130_fd_sc_hd__nor2_1
X_11258_ _15947_/Q _11268_/C _11202_/X vssd1 vssd1 vccd1 vccd1 _11258_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10209_ _10205_/Y _10216_/A _10208_/Y _10201_/C vssd1 vssd1 vccd1 vccd1 _10211_/B
+ sky130_fd_sc_hd__o211a_1
X_11189_ _15937_/Q _11197_/C _11188_/X vssd1 vssd1 vccd1 vccd1 _11189_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15997_ _16005_/CLK _15997_/D vssd1 vssd1 vccd1 vccd1 _15997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14948_ _14948_/A _14956_/B vssd1 vssd1 vccd1 vccd1 _14950_/A sky130_fd_sc_hd__or2_1
XFILLER_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14879_ _14879_/A vssd1 vssd1 vccd1 vccd1 _16465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16618_ input11/X _16618_/D vssd1 vssd1 vccd1 vccd1 _16618_/Q sky130_fd_sc_hd__dfxtp_1
X_16549_ _16551_/CLK _16549_/D vssd1 vssd1 vccd1 vccd1 _16549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09021_ _15541_/Q _09028_/C _08859_/X vssd1 vssd1 vccd1 vccd1 _09021_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09923_ _09921_/A _09921_/B _09920_/Y _09922_/Y vssd1 vssd1 vccd1 vccd1 _15718_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_131_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09854_ _09851_/X _09846_/B _09849_/B _09853_/Y vssd1 vssd1 vccd1 vccd1 _15703_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08805_ _09056_/A vssd1 vssd1 vccd1 vccd1 _08805_/X sky130_fd_sc_hd__clkbuf_4
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _09780_/Y _09783_/X _09784_/Y vssd1 vssd1 vccd1 vccd1 _15692_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08736_ _08870_/A _08736_/B vssd1 vssd1 vccd1 vccd1 _08736_/X sky130_fd_sc_hd__or2_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _08667_/A vssd1 vssd1 vccd1 vccd1 _08667_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _08854_/A vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10560_ _15837_/Q _10702_/B _10565_/C vssd1 vssd1 vccd1 vccd1 _10560_/Y sky130_fd_sc_hd__nand3_1
X_09219_ _15585_/Q _09220_/C _09364_/B vssd1 vssd1 vccd1 vccd1 _09222_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _10491_/A vssd1 vssd1 vccd1 vccd1 _15824_/D sky130_fd_sc_hd__clkbuf_1
X_12230_ _12230_/A _12230_/B _12234_/B vssd1 vssd1 vccd1 vccd1 _16083_/D sky130_fd_sc_hd__nor3_1
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ _12158_/Y _12159_/X _12160_/Y _12155_/C vssd1 vssd1 vccd1 vccd1 _12163_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11112_ _11266_/A vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__buf_2
XFILLER_150_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12092_ _16065_/Q _12100_/C _12036_/X vssd1 vssd1 vccd1 vccd1 _12092_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11043_ _11097_/A _11043_/B _11047_/B vssd1 vssd1 vccd1 vccd1 _15915_/D sky130_fd_sc_hd__nor3_1
X_15920_ _15365_/A _15920_/D vssd1 vssd1 vccd1 vccd1 _15920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15851_ _16595_/CLK _15851_/D vssd1 vssd1 vccd1 vccd1 _15851_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14802_ _14795_/C _14796_/C _14798_/Y _14800_/X vssd1 vssd1 vccd1 vccd1 _14803_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_36_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15782_ _15812_/CLK _15782_/D vssd1 vssd1 vccd1 vccd1 _15782_/Q sky130_fd_sc_hd__dfxtp_1
X_12994_ _16192_/Q _13001_/C _12879_/X vssd1 vssd1 vccd1 vccd1 _12997_/B sky130_fd_sc_hd__a21o_1
XFILLER_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14733_ _16444_/Q _14790_/B _14742_/C vssd1 vssd1 vccd1 vccd1 _14738_/A sky130_fd_sc_hd__and3_1
X_11945_ _16043_/Q _12060_/B _11950_/C vssd1 vssd1 vccd1 vccd1 _11945_/Y sky130_fd_sc_hd__nand3_1
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14664_ _14664_/A _14664_/B vssd1 vssd1 vccd1 vccd1 _14665_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11876_ _16034_/Q _11878_/C _11875_/X vssd1 vssd1 vccd1 vccd1 _11876_/Y sky130_fd_sc_hd__a21oi_1
X_16403_ _16607_/CLK _16403_/D vssd1 vssd1 vccd1 vccd1 _16403_/Q sky130_fd_sc_hd__dfxtp_1
X_13615_ _13615_/A vssd1 vssd1 vccd1 vccd1 _16279_/D sky130_fd_sc_hd__clkbuf_1
X_10827_ _11266_/A vssd1 vssd1 vccd1 vccd1 _10954_/A sky130_fd_sc_hd__buf_2
XFILLER_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14595_ _14595_/A vssd1 vssd1 vccd1 vccd1 _16420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16334_ _16346_/CLK _16334_/D vssd1 vssd1 vccd1 vccd1 _16334_/Q sky130_fd_sc_hd__dfxtp_2
X_13546_ _14669_/A vssd1 vssd1 vccd1 vccd1 _13546_/X sky130_fd_sc_hd__clkbuf_2
X_10758_ _10758_/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10759_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16265_ _16533_/Q _16265_/D vssd1 vssd1 vccd1 vccd1 _16265_/Q sky130_fd_sc_hd__dfxtp_1
X_13477_ _13498_/A _13477_/B _13481_/B vssd1 vssd1 vccd1 vccd1 _16259_/D sky130_fd_sc_hd__nor3_1
X_10689_ _10689_/A vssd1 vssd1 vccd1 vccd1 _15861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15216_ _15216_/A _15223_/B vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__or2_1
X_12428_ _16112_/Q _12435_/C _12316_/X vssd1 vssd1 vccd1 vccd1 _12431_/B sky130_fd_sc_hd__a21o_1
X_16196_ _16555_/Q _16196_/D vssd1 vssd1 vccd1 vccd1 _16196_/Q sky130_fd_sc_hd__dfxtp_1
X_15147_ _16511_/Q _15155_/C _10797_/B vssd1 vssd1 vccd1 vccd1 _15147_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ _12361_/B _12361_/C _12133_/X vssd1 vssd1 vccd1 vccd1 _12362_/B sky130_fd_sc_hd__o21ai_1
XFILLER_126_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15078_ _15079_/B _15079_/C _15079_/A vssd1 vssd1 vccd1 vccd1 _15080_/B sky130_fd_sc_hd__a21o_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14029_ _14308_/A vssd1 vssd1 vccd1 vccd1 _14029_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09570_ _09438_/X _09568_/B _09530_/X vssd1 vssd1 vccd1 vccd1 _09570_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08521_ _08521_/A _08521_/B vssd1 vssd1 vccd1 vccd1 _15307_/C sky130_fd_sc_hd__xor2_2
XFILLER_36_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08452_ _08504_/A _08504_/B vssd1 vssd1 vccd1 vccd1 _08505_/A sky130_fd_sc_hd__xnor2_2
XFILLER_91_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08383_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08455_/A sky130_fd_sc_hd__xnor2_2
XFILLER_149_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09004_ _08923_/X _09002_/A _08924_/X vssd1 vssd1 vccd1 vccd1 _09005_/B sky130_fd_sc_hd__o21ai_1
XFILLER_3_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09906_ _09946_/A _09906_/B _09910_/A vssd1 vssd1 vccd1 vccd1 _15715_/D sky130_fd_sc_hd__nor3_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09837_ _09837_/A vssd1 vssd1 vccd1 vccd1 _10308_/C sky130_fd_sc_hd__clkbuf_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09768_ _09768_/A vssd1 vssd1 vccd1 vccd1 _15689_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08730_/A _08719_/B _08723_/A vssd1 vssd1 vccd1 vccd1 _15472_/D sky130_fd_sc_hd__nor3_1
XFILLER_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09699_ _09699_/A vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _11730_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__or2_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _12225_/A vssd1 vssd1 vccd1 vccd1 _11891_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _16250_/Q _13623_/B _13401_/C vssd1 vssd1 vccd1 vccd1 _13400_/X sky130_fd_sc_hd__and3_1
X_10612_ _15848_/Q _10707_/B _10612_/C vssd1 vssd1 vccd1 vccd1 _10613_/B sky130_fd_sc_hd__and3_1
X_14380_ _16389_/Q _14486_/B _14380_/C vssd1 vssd1 vccd1 vccd1 _14389_/B sky130_fd_sc_hd__and3_1
X_11592_ _15994_/Q _11594_/C _11591_/X vssd1 vssd1 vccd1 vccd1 _11592_/Y sky130_fd_sc_hd__a21oi_1
X_13331_ _13332_/B _13332_/C _13332_/A vssd1 vssd1 vccd1 vccd1 _13333_/B sky130_fd_sc_hd__a21o_1
X_10543_ _10543_/A vssd1 vssd1 vccd1 vccd1 _15833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16050_ _16118_/CLK _16050_/D vssd1 vssd1 vccd1 vccd1 _16050_/Q sky130_fd_sc_hd__dfxtp_1
X_13262_ _13260_/A _13260_/B _13261_/X vssd1 vssd1 vccd1 vccd1 _16228_/D sky130_fd_sc_hd__a21oi_1
X_10474_ _10418_/X _10471_/B _10473_/X vssd1 vssd1 vccd1 vccd1 _10474_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_142_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15001_ _16486_/Q _15055_/B _15001_/C vssd1 vssd1 vccd1 vccd1 _15009_/B sky130_fd_sc_hd__and3_1
X_12213_ _12209_/Y _12210_/X _12212_/Y _12207_/C vssd1 vssd1 vccd1 vccd1 _12215_/B
+ sky130_fd_sc_hd__o211ai_1
X_13193_ _16220_/Q _13305_/B _13193_/C vssd1 vssd1 vccd1 vccd1 _13201_/A sky130_fd_sc_hd__and3_1
XFILLER_2_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12144_ _12230_/A _12144_/B _12148_/A vssd1 vssd1 vccd1 vccd1 _16070_/D sky130_fd_sc_hd__nor3_1
XFILLER_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16658__63 vssd1 vssd1 vccd1 vccd1 _16658__63/HI _16734_/A sky130_fd_sc_hd__conb_1
X_12075_ _12113_/A _12075_/B _12075_/C vssd1 vssd1 vccd1 vccd1 _12076_/A sky130_fd_sc_hd__and3_1
XFILLER_2_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11026_ _15913_/Q _11026_/B _11026_/C vssd1 vssd1 vccd1 vccd1 _11026_/Y sky130_fd_sc_hd__nand3_1
X_15903_ _16553_/Q _15903_/D vssd1 vssd1 vccd1 vccd1 _15903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15834_ _16595_/CLK _15834_/D vssd1 vssd1 vccd1 vccd1 _15834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15765_ _15812_/CLK _15765_/D vssd1 vssd1 vccd1 vccd1 _15765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12977_ _12977_/A _12977_/B vssd1 vssd1 vccd1 vccd1 _12978_/B sky130_fd_sc_hd__nor2_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14716_ _16441_/Q _14770_/B _14716_/C vssd1 vssd1 vccd1 vccd1 _14724_/B sky130_fd_sc_hd__and3_1
X_11928_ _16042_/Q _11928_/B _11930_/C vssd1 vssd1 vccd1 vccd1 _11928_/X sky130_fd_sc_hd__and3_1
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15696_ _15791_/CLK _15696_/D vssd1 vssd1 vccd1 vccd1 _15696_/Q sky130_fd_sc_hd__dfxtp_4
X_14647_ _14647_/A vssd1 vssd1 vccd1 vccd1 _14875_/B sky130_fd_sc_hd__clkbuf_2
X_11859_ _16031_/Q _11897_/C _11802_/X vssd1 vssd1 vccd1 vccd1 _11861_/B sky130_fd_sc_hd__a21oi_1
XFILLER_20_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_18 _14790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 _09849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ _14571_/C _14572_/C _14575_/Y _14576_/X vssd1 vssd1 vccd1 vccd1 _14579_/C
+ sky130_fd_sc_hd__a211o_1
X_16317_ _16389_/CLK _16317_/D vssd1 vssd1 vccd1 vccd1 _16317_/Q sky130_fd_sc_hd__dfxtp_1
X_13529_ _14092_/A vssd1 vssd1 vccd1 vccd1 _13643_/A sky130_fd_sc_hd__buf_2
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16248_ _16261_/CLK _16248_/D vssd1 vssd1 vccd1 vccd1 _16248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16179_ _16237_/CLK _16179_/D vssd1 vssd1 vccd1 vccd1 _16179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07952_ _16556_/Q vssd1 vssd1 vccd1 vccd1 _10767_/A sky130_fd_sc_hd__inv_2
XFILLER_102_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07883_ _16597_/Q vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__clkinv_2
XFILLER_68_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09622_ _09625_/C vssd1 vssd1 vccd1 vccd1 _09636_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09553_ _09595_/A _09553_/B _09556_/B vssd1 vssd1 vccd1 vccd1 _15645_/D sky130_fd_sc_hd__nor3_1
XFILLER_36_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08504_ _08504_/A _08504_/B vssd1 vssd1 vccd1 vccd1 _08509_/A sky130_fd_sc_hd__or2_1
XFILLER_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09484_ _09299_/X _09481_/B _09483_/Y vssd1 vssd1 vccd1 vccd1 _15631_/D sky130_fd_sc_hd__o21a_1
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ _08435_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08435_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08366_ _08366_/A _08366_/B vssd1 vssd1 vccd1 vccd1 _08437_/A sky130_fd_sc_hd__xnor2_2
XFILLER_149_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08297_ _09178_/C _07900_/B _08296_/X vssd1 vssd1 vccd1 vccd1 _08299_/A sky130_fd_sc_hd__o21ai_1
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10190_ _15773_/Q _10190_/B _10190_/C vssd1 vssd1 vccd1 vccd1 _10190_/X sky130_fd_sc_hd__and3_1
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12900_ _12900_/A vssd1 vssd1 vccd1 vccd1 _16177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13880_ _13878_/A _13878_/B _13879_/X vssd1 vssd1 vccd1 vccd1 _16316_/D sky130_fd_sc_hd__a21oi_1
XFILLER_46_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _12847_/A _12831_/B _12831_/C vssd1 vssd1 vccd1 vccd1 _12832_/A sky130_fd_sc_hd__and3_1
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15550_ _16551_/CLK _15550_/D vssd1 vssd1 vccd1 vccd1 _15550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12796_/A _12762_/B _12766_/A vssd1 vssd1 vccd1 vccd1 _16158_/D sky130_fd_sc_hd__nor3_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _16424_/Q vssd1 vssd1 vccd1 vccd1 _14516_/C sky130_fd_sc_hd__inv_2
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11713_ _16011_/Q _11936_/B _11721_/C vssd1 vssd1 vccd1 vccd1 _11713_/X sky130_fd_sc_hd__and3_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _16570_/CLK _15481_/D vssd1 vssd1 vccd1 vccd1 _15481_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12693_ _12693_/A _12701_/B vssd1 vssd1 vccd1 vccd1 _12695_/A sky130_fd_sc_hd__or2_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _16397_/Q _14433_/C _14265_/X vssd1 vssd1 vccd1 vccd1 _14434_/A sky130_fd_sc_hd__a21oi_1
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11644_ _16002_/Q _11644_/B _11648_/C vssd1 vssd1 vccd1 vccd1 _11644_/X sky130_fd_sc_hd__and3_1
X_14363_ _16387_/Q _14373_/C _14308_/X vssd1 vssd1 vccd1 vccd1 _14363_/Y sky130_fd_sc_hd__a21oi_1
X_11575_ _11607_/C vssd1 vssd1 vccd1 vccd1 _11613_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16102_ _16118_/CLK _16102_/D vssd1 vssd1 vccd1 vccd1 _16102_/Q sky130_fd_sc_hd__dfxtp_2
X_13314_ _13314_/A _13314_/B vssd1 vssd1 vccd1 vccd1 _13319_/C sky130_fd_sc_hd__nor2_1
XFILLER_128_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10526_ _10526_/A vssd1 vssd1 vccd1 vccd1 _10526_/X sky130_fd_sc_hd__clkbuf_2
X_14294_ _14858_/A vssd1 vssd1 vccd1 vccd1 _14294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16033_ _16118_/CLK _16033_/D vssd1 vssd1 vccd1 vccd1 _16033_/Q sky130_fd_sc_hd__dfxtp_1
X_13245_ _13243_/Y _13238_/C _13240_/Y _13241_/X vssd1 vssd1 vccd1 vccd1 _13246_/C
+ sky130_fd_sc_hd__a211o_1
X_10457_ _15820_/Q _10652_/B _10457_/C vssd1 vssd1 vccd1 vccd1 _10465_/A sky130_fd_sc_hd__and3_1
XFILLER_108_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13176_ _16218_/Q _13178_/C _13006_/X vssd1 vssd1 vccd1 vccd1 _13176_/Y sky130_fd_sc_hd__a21oi_1
X_10388_ _15809_/Q _10494_/B _10388_/C vssd1 vssd1 vccd1 vccd1 _10388_/X sky130_fd_sc_hd__and3_1
XFILLER_124_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ _12127_/A _12127_/B vssd1 vssd1 vccd1 vccd1 _12128_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12058_ _16060_/Q _12065_/C _12000_/X vssd1 vssd1 vccd1 vccd1 _12058_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11009_ _15911_/Q _11118_/B _11018_/C vssd1 vssd1 vccd1 vccd1 _11014_/A sky130_fd_sc_hd__and3_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15817_ _16570_/CLK _15817_/D vssd1 vssd1 vccd1 vccd1 _15817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15748_ _15812_/CLK _15748_/D vssd1 vssd1 vccd1 vccd1 _15748_/Q sky130_fd_sc_hd__dfxtp_1
X_15679_ _15791_/CLK _15679_/D vssd1 vssd1 vccd1 vccd1 _15679_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08220_ _08220_/A _08220_/B vssd1 vssd1 vccd1 vccd1 _08454_/B sky130_fd_sc_hd__xnor2_4
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08151_ _13212_/A _08151_/B vssd1 vssd1 vccd1 vccd1 _08151_/X sky130_fd_sc_hd__or2_1
XFILLER_119_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08082_ _08082_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08083_/B sky130_fd_sc_hd__nand2_2
XFILLER_106_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08984_ _09998_/B vssd1 vssd1 vccd1 vccd1 _09145_/B sky130_fd_sc_hd__clkbuf_2
X_07935_ _16605_/Q vssd1 vssd1 vccd1 vccd1 _13551_/A sky130_fd_sc_hd__clkinv_2
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07866_ _15822_/Q vssd1 vssd1 vccd1 vccd1 _10379_/C sky130_fd_sc_hd__inv_2
XFILLER_29_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09605_ _15659_/Q _09603_/C _09604_/X vssd1 vssd1 vccd1 vccd1 _09606_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07797_ _07799_/A vssd1 vssd1 vccd1 vccd1 _07797_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09536_ _09756_/A vssd1 vssd1 vccd1 vccd1 _09536_/X sky130_fd_sc_hd__buf_2
XFILLER_43_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09467_ _09467_/A _09467_/B vssd1 vssd1 vccd1 vccd1 _09467_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ _15291_/A _08418_/B vssd1 vssd1 vccd1 vccd1 _08419_/B sky130_fd_sc_hd__nand2_1
X_09398_ _09398_/A _09398_/B vssd1 vssd1 vccd1 vccd1 _15614_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08349_ _08226_/A _08226_/B _08348_/X vssd1 vssd1 vccd1 vccd1 _08366_/A sky130_fd_sc_hd__a21bo_1
XFILLER_137_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _11360_/A vssd1 vssd1 vccd1 vccd1 _11594_/B sky130_fd_sc_hd__buf_2
XFILLER_138_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10311_ _10311_/A _10311_/B _10315_/B vssd1 vssd1 vccd1 vccd1 _15791_/D sky130_fd_sc_hd__nor3_1
XFILLER_3_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11291_ _15951_/Q _11328_/C _11233_/X vssd1 vssd1 vccd1 vccd1 _11293_/B sky130_fd_sc_hd__a21oi_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13030_ _13030_/A _13030_/B vssd1 vssd1 vccd1 vccd1 _13031_/B sky130_fd_sc_hd__nor2_1
X_10242_ _10242_/A vssd1 vssd1 vccd1 vccd1 _15779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10173_ _10190_/C vssd1 vssd1 vccd1 vccd1 _10206_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16628__33 vssd1 vssd1 vccd1 vccd1 _16628__33/HI _16694_/A sky130_fd_sc_hd__conb_1
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14981_ _16483_/Q _15033_/B _14982_/C vssd1 vssd1 vccd1 vccd1 _14981_/X sky130_fd_sc_hd__and3_1
XFILLER_75_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16720_ _16720_/A _07824_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13932_ _14210_/A vssd1 vssd1 vccd1 vccd1 _14158_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13863_ _16314_/Q _14032_/B _13869_/C vssd1 vssd1 vccd1 vccd1 _13863_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15602_ _16551_/CLK _15602_/D vssd1 vssd1 vccd1 vccd1 _15602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12814_ _12828_/C vssd1 vssd1 vccd1 vccd1 _12836_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13794_ _13792_/Y _13793_/X _13789_/C _13790_/C vssd1 vssd1 vccd1 vccd1 _13796_/B
+ sky130_fd_sc_hd__o211ai_1
X_16582_ _16595_/CLK _16582_/D vssd1 vssd1 vccd1 vccd1 _16582_/Q sky130_fd_sc_hd__dfxtp_1
X_15533_ _16551_/CLK _15533_/D vssd1 vssd1 vccd1 vccd1 _15533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _16157_/Q _12798_/B _12745_/C vssd1 vssd1 vccd1 vccd1 _12753_/B sky130_fd_sc_hd__and3_1
XFILLER_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15464_ _16570_/CLK _15464_/D vssd1 vssd1 vccd1 vccd1 _15464_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _16147_/Q _12784_/B _12685_/C vssd1 vssd1 vccd1 vccd1 _12676_/X sky130_fd_sc_hd__and3_1
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ _14412_/Y _14413_/X _14414_/Y _14409_/C vssd1 vssd1 vccd1 vccd1 _14417_/B
+ sky130_fd_sc_hd__o211ai_1
X_11627_ _11662_/C vssd1 vssd1 vccd1 vccd1 _11668_/C sky130_fd_sc_hd__clkbuf_2
X_15395_ _16061_/Q _16060_/Q _16059_/Q _15391_/X vssd1 vssd1 vccd1 vccd1 _16578_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_129_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14346_ _14347_/B _14347_/C _14347_/A vssd1 vssd1 vccd1 vccd1 _14348_/B sky130_fd_sc_hd__a21o_1
X_11558_ _11666_/A _11558_/B _11562_/B vssd1 vssd1 vccd1 vccd1 _15987_/D sky130_fd_sc_hd__nor3_1
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _15829_/Q _10652_/B _10509_/C vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__and3_1
XFILLER_128_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14277_ _14314_/A _14277_/B _14277_/C vssd1 vssd1 vccd1 vccd1 _14278_/A sky130_fd_sc_hd__and3_1
X_11489_ _11486_/Y _11487_/X _11488_/Y _11483_/C vssd1 vssd1 vccd1 vccd1 _11491_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_143_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16016_ _16554_/Q _16016_/D vssd1 vssd1 vccd1 vccd1 _16016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13228_ _16225_/Q _13336_/B _13228_/C vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__and3_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13725_/A vssd1 vssd1 vccd1 vccd1 _13383_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ _09374_/A _09321_/B _09325_/A vssd1 vssd1 vccd1 vccd1 _15598_/D sky130_fd_sc_hd__nor3_1
X_09252_ _09943_/A vssd1 vssd1 vccd1 vccd1 _09252_/X sky130_fd_sc_hd__buf_2
XFILLER_139_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08203_ _08204_/A _08204_/B _08204_/C vssd1 vssd1 vccd1 vccd1 _08357_/A sky130_fd_sc_hd__a21oi_2
XFILLER_138_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ _15577_/Q _09192_/C _09063_/X vssd1 vssd1 vccd1 vccd1 _09183_/Y sky130_fd_sc_hd__a21oi_1
X_08134_ _08332_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08135_/B sky130_fd_sc_hd__xnor2_2
XFILLER_135_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08065_ _09496_/C _08065_/B vssd1 vssd1 vccd1 vccd1 _08066_/B sky130_fd_sc_hd__xnor2_4
XFILLER_134_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08967_ _08883_/X _08965_/A _08966_/Y vssd1 vssd1 vccd1 vccd1 _15524_/D sky130_fd_sc_hd__o21a_1
XFILLER_103_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07918_ _15858_/Q vssd1 vssd1 vccd1 vccd1 _10583_/C sky130_fd_sc_hd__clkinv_2
XFILLER_69_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08898_ _08898_/A _08898_/B _08898_/C vssd1 vssd1 vccd1 vccd1 _08899_/C sky130_fd_sc_hd__nand3_1
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07849_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07849_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _15891_/Q _11084_/B _10868_/C vssd1 vssd1 vccd1 vccd1 _10860_/X sky130_fd_sc_hd__and3_1
XFILLER_25_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ _15641_/Q _09692_/B _09519_/C vssd1 vssd1 vccd1 vccd1 _09519_/X sky130_fd_sc_hd__and3_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _15880_/Q _11026_/B _10791_/C vssd1 vssd1 vccd1 vccd1 _10791_/Y sky130_fd_sc_hd__nand3_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _16587_/Q vssd1 vssd1 vccd1 vccd1 _12545_/C sky130_fd_sc_hd__inv_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _16117_/Q _12462_/C _12292_/X vssd1 vssd1 vccd1 vccd1 _12463_/A sky130_fd_sc_hd__a21oi_1
XFILLER_149_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14200_ _15048_/A vssd1 vssd1 vccd1 vccd1 _14427_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_11412_ _15969_/Q _11638_/B _11412_/C vssd1 vssd1 vccd1 vccd1 _11412_/X sky130_fd_sc_hd__and3_1
X_15180_ _15180_/A _15180_/B _15184_/A vssd1 vssd1 vccd1 vccd1 _16515_/D sky130_fd_sc_hd__nor3_1
XFILLER_137_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12392_ _16107_/Q _12402_/C _12337_/X vssd1 vssd1 vccd1 vccd1 _12392_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _14131_/A vssd1 vssd1 vccd1 vccd1 _16352_/D sky130_fd_sc_hd__clkbuf_1
X_11343_ _15959_/Q _11381_/C _11233_/X vssd1 vssd1 vccd1 vccd1 _11345_/B sky130_fd_sc_hd__a21oi_1
XFILLER_126_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14062_ _16343_/Q _14227_/B _14072_/C vssd1 vssd1 vccd1 vccd1 _14068_/A sky130_fd_sc_hd__and3_1
X_11274_ _15949_/Q _11275_/C _11158_/X vssd1 vssd1 vccd1 vccd1 _11276_/A sky130_fd_sc_hd__a21oi_1
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13013_ _13013_/A vssd1 vssd1 vccd1 vccd1 _16193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10225_ _10168_/X _10222_/B _10224_/X vssd1 vssd1 vccd1 vccd1 _10225_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10156_ _10179_/A _10156_/B _10160_/B vssd1 vssd1 vccd1 vccd1 _15764_/D sky130_fd_sc_hd__nor3_1
XFILLER_66_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10087_ _10085_/Y _10086_/X _10081_/C _10082_/C vssd1 vssd1 vccd1 vccd1 _10089_/B
+ sky130_fd_sc_hd__o211ai_1
X_14964_ _16480_/Q _15001_/C _14906_/X vssd1 vssd1 vccd1 vccd1 _14966_/B sky130_fd_sc_hd__a21oi_1
X_16703_ _16703_/A _07803_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
X_13915_ _16322_/Q _14032_/B _13923_/C vssd1 vssd1 vccd1 vccd1 _13915_/Y sky130_fd_sc_hd__nand3_1
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14895_ _14895_/A vssd1 vssd1 vccd1 vccd1 _15117_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13846_ _13846_/A vssd1 vssd1 vccd1 vccd1 _16311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16565_ _16570_/CLK _16565_/D vssd1 vssd1 vccd1 vccd1 _16565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13777_ _13777_/A vssd1 vssd1 vccd1 vccd1 _13793_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10989_ _10987_/Y _10981_/C _10984_/Y _10994_/A vssd1 vssd1 vccd1 vccd1 _10994_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15516_ _16551_/CLK _15516_/D vssd1 vssd1 vccd1 vccd1 _15516_/Q sky130_fd_sc_hd__dfxtp_1
X_12728_ _12726_/Y _12721_/C _12724_/Y _12725_/X vssd1 vssd1 vccd1 vccd1 _12729_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16496_ _16607_/CLK _16496_/D vssd1 vssd1 vccd1 vccd1 _16496_/Q sky130_fd_sc_hd__dfxtp_1
X_12659_ _12659_/A _12659_/B _12659_/C vssd1 vssd1 vccd1 vccd1 _12660_/C sky130_fd_sc_hd__nand3_1
X_15447_ _16570_/CLK _15447_/D vssd1 vssd1 vccd1 vccd1 _15447_/Q sky130_fd_sc_hd__dfxtp_1
X_15378_ _15378_/A vssd1 vssd1 vccd1 vccd1 _15378_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ _14439_/A vssd1 vssd1 vccd1 vccd1 _14369_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _09951_/A _09870_/B _09870_/C vssd1 vssd1 vccd1 vccd1 _09871_/A sky130_fd_sc_hd__and3_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _10393_/A vssd1 vssd1 vccd1 vccd1 _08991_/B sky130_fd_sc_hd__clkbuf_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08921_/A _08921_/B _08752_/C vssd1 vssd1 vccd1 vccd1 _08754_/A sky130_fd_sc_hd__and3_1
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08683_ _15469_/Q _08689_/C _08604_/X vssd1 vssd1 vccd1 vccd1 _08683_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09304_ _09750_/A vssd1 vssd1 vccd1 vccd1 _09304_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ _09849_/A _09235_/B vssd1 vssd1 vccd1 vccd1 _09235_/X sky130_fd_sc_hd__or2_1
XFILLER_22_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09166_ _09125_/X _09162_/A _09126_/X vssd1 vssd1 vccd1 vccd1 _09167_/B sky130_fd_sc_hd__o21ai_1
XFILLER_119_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08117_ _11339_/A _07898_/B _08116_/X vssd1 vssd1 vccd1 vccd1 _08145_/A sky130_fd_sc_hd__o21ai_1
XFILLER_108_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09097_ _09148_/A _09097_/B _09101_/A vssd1 vssd1 vccd1 vccd1 _15553_/D sky130_fd_sc_hd__nor3_1
XFILLER_135_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08048_ _14675_/A _08048_/B vssd1 vssd1 vccd1 vccd1 _08239_/B sky130_fd_sc_hd__xnor2_2
XFILLER_150_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10010_ _15740_/Q _10009_/C _08629_/A vssd1 vssd1 vccd1 vccd1 _10011_/B sky130_fd_sc_hd__a21o_1
XFILLER_88_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09999_ _09997_/Y _10004_/A _09994_/C _09995_/C vssd1 vssd1 vccd1 vccd1 _10001_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11961_ _11998_/A _11961_/B _11961_/C vssd1 vssd1 vccd1 vccd1 _11962_/A sky130_fd_sc_hd__and3_1
XFILLER_72_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10912_ _15898_/Q _10914_/C _14932_/A vssd1 vssd1 vccd1 vccd1 _10912_/Y sky130_fd_sc_hd__a21oi_1
X_13700_ _16292_/Q _13869_/B _13700_/C vssd1 vssd1 vccd1 vccd1 _13711_/A sky130_fd_sc_hd__and3_1
XFILLER_45_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14680_ _16435_/Q _14790_/B _14689_/C vssd1 vssd1 vccd1 vccd1 _14685_/A sky130_fd_sc_hd__and3_1
XFILLER_71_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11892_ _16035_/Q _12060_/B _11897_/C vssd1 vssd1 vccd1 vccd1 _11892_/Y sky130_fd_sc_hd__nand3_1
XFILLER_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13631_ _16283_/Q _13631_/B _13639_/C vssd1 vssd1 vccd1 vccd1 _13631_/X sky130_fd_sc_hd__and3_1
X_10843_ _11978_/A vssd1 vssd1 vccd1 vccd1 _11070_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13562_ _13583_/A _13562_/B _13562_/C vssd1 vssd1 vccd1 vccd1 _13563_/A sky130_fd_sc_hd__and3_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16350_ _16389_/CLK _16350_/D vssd1 vssd1 vccd1 vccd1 _16350_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10774_ _15879_/Q _10782_/C _15235_/B vssd1 vssd1 vccd1 vccd1 _10777_/B sky130_fd_sc_hd__a21o_1
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15301_ _15301_/A _15301_/B vssd1 vssd1 vccd1 vccd1 _15303_/A sky130_fd_sc_hd__nand2_1
X_12513_ _12511_/Y _12505_/C _12507_/Y _12518_/A vssd1 vssd1 vccd1 vccd1 _12518_/B
+ sky130_fd_sc_hd__a211oi_1
X_16281_ _16533_/Q _16281_/D vssd1 vssd1 vccd1 vccd1 _16281_/Q sky130_fd_sc_hd__dfxtp_1
X_13493_ _13514_/C vssd1 vssd1 vccd1 vccd1 _13531_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15232_ _16525_/Q _15232_/B _15241_/C vssd1 vssd1 vccd1 vccd1 _15237_/A sky130_fd_sc_hd__and3_1
X_12444_ _12441_/Y _12442_/X _12443_/Y _12438_/C vssd1 vssd1 vccd1 vccd1 _12446_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ _15163_/A _15163_/B vssd1 vssd1 vccd1 vccd1 _15164_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12375_ _12376_/B _12376_/C _12376_/A vssd1 vssd1 vccd1 vccd1 _12377_/B sky130_fd_sc_hd__a21o_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14114_ _14127_/C vssd1 vssd1 vccd1 vccd1 _14135_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11326_ _11379_/A _11326_/B _11330_/B vssd1 vssd1 vccd1 vccd1 _15955_/D sky130_fd_sc_hd__nor3_1
X_15094_ _15094_/A vssd1 vssd1 vccd1 vccd1 _16500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14045_ _14045_/A _14053_/B vssd1 vssd1 vccd1 vccd1 _14047_/A sky130_fd_sc_hd__or2_1
X_11257_ _11257_/A vssd1 vssd1 vccd1 vccd1 _15945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10208_ _15774_/Q _10458_/B _10214_/C vssd1 vssd1 vccd1 vccd1 _10208_/Y sky130_fd_sc_hd__nand3_1
XFILLER_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11188_ _13060_/A vssd1 vssd1 vccd1 vccd1 _11188_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10139_ _15765_/Q _10152_/C _10138_/X vssd1 vssd1 vccd1 vccd1 _10139_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15996_ _16005_/CLK _15996_/D vssd1 vssd1 vccd1 vccd1 _15996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14947_ _16477_/Q _15055_/B _14947_/C vssd1 vssd1 vccd1 vccd1 _14956_/B sky130_fd_sc_hd__and3_1
XFILLER_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14878_ _14878_/A _14878_/B _14878_/C vssd1 vssd1 vccd1 vccd1 _14879_/A sky130_fd_sc_hd__and3_1
XFILLER_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16617_ input11/X _16617_/D vssd1 vssd1 vccd1 vccd1 _16617_/Q sky130_fd_sc_hd__dfxtp_1
X_13829_ _14669_/A vssd1 vssd1 vccd1 vccd1 _13829_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16548_ _16551_/CLK _16548_/D vssd1 vssd1 vccd1 vccd1 _16548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16479_ _16607_/CLK _16479_/D vssd1 vssd1 vccd1 vccd1 _16479_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ _09020_/A vssd1 vssd1 vccd1 vccd1 _15536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09922_ _09921_/X _09920_/Y _08700_/A vssd1 vssd1 vccd1 vccd1 _09922_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09853_ _10065_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09853_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _08846_/A _08804_/B _08809_/A vssd1 vssd1 vccd1 vccd1 _15490_/D sky130_fd_sc_hd__nor3_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09784_ _09780_/Y _09783_/X _09750_/X vssd1 vssd1 vccd1 vccd1 _09784_/Y sky130_fd_sc_hd__a21oi_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _08735_/A _08735_/B vssd1 vssd1 vccd1 vccd1 _08736_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _09126_/A vssd1 vssd1 vccd1 vccd1 _08667_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08597_ _10060_/A vssd1 vssd1 vccd1 vccd1 _08854_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09218_ _09629_/A vssd1 vssd1 vccd1 vccd1 _09364_/B sky130_fd_sc_hd__buf_2
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10490_ _10497_/A _10490_/B _10490_/C vssd1 vssd1 vccd1 vccd1 _10491_/A sky130_fd_sc_hd__and3_1
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09149_ _15569_/Q _09150_/C _08989_/X vssd1 vssd1 vccd1 vccd1 _09151_/A sky130_fd_sc_hd__a21oi_1
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12160_ _16073_/Q _12160_/B _12160_/C vssd1 vssd1 vccd1 vccd1 _12160_/Y sky130_fd_sc_hd__nand3_1
XFILLER_107_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11111_ _11111_/A vssd1 vssd1 vccd1 vccd1 _15925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12091_ _12091_/A vssd1 vssd1 vccd1 vccd1 _16063_/D sky130_fd_sc_hd__clkbuf_1
X_11042_ _11040_/Y _11036_/C _11038_/Y _11047_/A vssd1 vssd1 vccd1 vccd1 _11047_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_104_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15850_ _16595_/CLK _15850_/D vssd1 vssd1 vccd1 vccd1 _15850_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14801_ _14798_/Y _14800_/X _14795_/C _14796_/C vssd1 vssd1 vccd1 vccd1 _14803_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15781_ _15812_/CLK _15781_/D vssd1 vssd1 vccd1 vccd1 _15781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12993_ _13080_/A _12993_/B _12997_/A vssd1 vssd1 vccd1 vccd1 _16190_/D sky130_fd_sc_hd__nor3_1
X_14732_ _16444_/Q _14770_/C _14621_/X vssd1 vssd1 vccd1 vccd1 _14734_/B sky130_fd_sc_hd__a21oi_1
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11944_ _16044_/Q _12173_/B _11944_/C vssd1 vssd1 vccd1 vccd1 _11952_/A sky130_fd_sc_hd__and3_1
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14663_ _14663_/A _14671_/B vssd1 vssd1 vccd1 vccd1 _14665_/A sky130_fd_sc_hd__or2_1
X_11875_ _13006_/A vssd1 vssd1 vccd1 vccd1 _11875_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16402_ _16607_/CLK _16402_/D vssd1 vssd1 vccd1 vccd1 _16402_/Q sky130_fd_sc_hd__dfxtp_1
X_13614_ _13635_/A _13614_/B _13614_/C vssd1 vssd1 vccd1 vccd1 _13615_/A sky130_fd_sc_hd__and3_1
XFILLER_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10826_ _15875_/Q _15874_/Q _15873_/Q _10719_/X vssd1 vssd1 vccd1 vccd1 _15885_/D
+ sky130_fd_sc_hd__o31a_1
X_14594_ _14594_/A _14594_/B _14594_/C vssd1 vssd1 vccd1 vccd1 _14595_/A sky130_fd_sc_hd__and3_1
X_16333_ _16346_/CLK _16333_/D vssd1 vssd1 vccd1 vccd1 _16333_/Q sky130_fd_sc_hd__dfxtp_1
X_10757_ _10757_/A _10757_/B vssd1 vssd1 vccd1 vccd1 _10758_/B sky130_fd_sc_hd__nor2_1
X_13545_ _13545_/A vssd1 vssd1 vccd1 vccd1 _14669_/A sky130_fd_sc_hd__buf_4
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16264_ _16533_/Q _16264_/D vssd1 vssd1 vccd1 vccd1 _16264_/Q sky130_fd_sc_hd__dfxtp_1
X_13476_ _13474_/Y _13470_/C _13472_/Y _13481_/A vssd1 vssd1 vccd1 vccd1 _13481_/B
+ sky130_fd_sc_hd__a211oi_1
X_10688_ _10738_/A _10688_/B _10688_/C vssd1 vssd1 vccd1 vccd1 _10689_/A sky130_fd_sc_hd__and3_1
XFILLER_145_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15215_ _16522_/Q _15267_/B _15215_/C vssd1 vssd1 vccd1 vccd1 _15223_/B sky130_fd_sc_hd__and3_1
X_12427_ _12514_/A _12427_/B _12431_/A vssd1 vssd1 vccd1 vccd1 _16110_/D sky130_fd_sc_hd__nor3_1
X_16195_ _16555_/Q _16195_/D vssd1 vssd1 vccd1 vccd1 _16195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15146_ _15146_/A vssd1 vssd1 vccd1 vccd1 _16509_/D sky130_fd_sc_hd__clkbuf_1
X_12358_ _12468_/A vssd1 vssd1 vccd1 vccd1 _12398_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11309_ _15953_/Q _11309_/B _11309_/C vssd1 vssd1 vccd1 vccd1 _11309_/Y sky130_fd_sc_hd__nand3_1
XFILLER_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15077_ _16499_/Q _15129_/B _15083_/C vssd1 vssd1 vccd1 vccd1 _15079_/C sky130_fd_sc_hd__nand3_1
X_12289_ _12286_/Y _12298_/A _12288_/Y _12283_/C vssd1 vssd1 vccd1 vccd1 _12291_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14028_ _14028_/A vssd1 vssd1 vccd1 vccd1 _16337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15979_ _16005_/CLK _15979_/D vssd1 vssd1 vccd1 vccd1 _15979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08520_ _08414_/A _08414_/B _08480_/A _08519_/X vssd1 vssd1 vccd1 vccd1 _08521_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08451_ _08357_/A _08357_/B _08450_/Y vssd1 vssd1 vccd1 vccd1 _08504_/B sky130_fd_sc_hd__a21oi_2
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08382_ _08253_/A _08252_/B _08252_/A vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__o21ba_1
XFILLER_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09003_ _09124_/A _09124_/B _09003_/C vssd1 vssd1 vccd1 vccd1 _09005_/A sky130_fd_sc_hd__and3_1
XFILLER_117_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09905_ _15718_/Q _09945_/B _09905_/C vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__and3_1
X_09836_ _15703_/Q _10307_/C _09836_/C vssd1 vssd1 vccd1 vccd1 _09847_/A sky130_fd_sc_hd__and3_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _09810_/A _09767_/B _09767_/C vssd1 vssd1 vccd1 vccd1 _09768_/A sky130_fd_sc_hd__and3_1
XFILLER_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _15476_/Q _08845_/B _08721_/C vssd1 vssd1 vccd1 vccd1 _08723_/A sky130_fd_sc_hd__and3_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09698_ _09698_/A vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _14828_/A vssd1 vssd1 vccd1 vccd1 _09164_/A sky130_fd_sc_hd__clkbuf_8
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _16004_/Q _11668_/C _11434_/X vssd1 vssd1 vccd1 vccd1 _11660_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _15848_/Q _10612_/C _08748_/A vssd1 vssd1 vccd1 vccd1 _10613_/A sky130_fd_sc_hd__a21oi_1
X_11591_ _13521_/A vssd1 vssd1 vccd1 vccd1 _11591_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13330_ _16240_/Q _13445_/B _13336_/C vssd1 vssd1 vccd1 vccd1 _13332_/C sky130_fd_sc_hd__nand3_1
XFILLER_10_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10542_ _10589_/A _10542_/B _10542_/C vssd1 vssd1 vccd1 vccd1 _10543_/A sky130_fd_sc_hd__and3_1
XFILLER_127_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _13315_/A _13266_/C vssd1 vssd1 vccd1 vccd1 _13261_/X sky130_fd_sc_hd__or2_1
XFILLER_10_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10473_ _10716_/A vssd1 vssd1 vccd1 vccd1 _10473_/X sky130_fd_sc_hd__clkbuf_2
X_15000_ _16486_/Q _15001_/C _14828_/X vssd1 vssd1 vccd1 vccd1 _15002_/A sky130_fd_sc_hd__a21oi_1
X_12212_ _16081_/Q _12443_/B _12212_/C vssd1 vssd1 vccd1 vccd1 _12212_/Y sky130_fd_sc_hd__nand3_1
XFILLER_136_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ _16220_/Q _13199_/C _13133_/X vssd1 vssd1 vccd1 vccd1 _13192_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12143_ _16071_/Q _12252_/B _12152_/C vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__and3_1
XFILLER_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12074_ _12304_/A _12074_/B _12074_/C vssd1 vssd1 vccd1 vccd1 _12075_/C sky130_fd_sc_hd__or3_1
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11025_ _15914_/Q _11076_/B _11026_/C vssd1 vssd1 vccd1 vccd1 _11025_/X sky130_fd_sc_hd__and3_1
X_15902_ _16553_/Q _15902_/D vssd1 vssd1 vccd1 vccd1 _15902_/Q sky130_fd_sc_hd__dfxtp_2
X_15833_ _16595_/CLK _15833_/D vssd1 vssd1 vccd1 vccd1 _15833_/Q sky130_fd_sc_hd__dfxtp_2
X_16673__78 vssd1 vssd1 vccd1 vccd1 _16673__78/HI _16749_/A sky130_fd_sc_hd__conb_1
XFILLER_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15764_ _15791_/CLK _15764_/D vssd1 vssd1 vccd1 vccd1 _15764_/Q sky130_fd_sc_hd__dfxtp_1
X_12976_ _12976_/A _12984_/B vssd1 vssd1 vccd1 vccd1 _12978_/A sky130_fd_sc_hd__or2_1
XFILLER_18_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14715_ _16441_/Q _14716_/C _14544_/X vssd1 vssd1 vccd1 vccd1 _14717_/A sky130_fd_sc_hd__a21oi_1
X_11927_ _16042_/Q _11930_/C _11875_/X vssd1 vssd1 vccd1 vccd1 _11927_/Y sky130_fd_sc_hd__a21oi_1
X_15695_ _15791_/CLK _15695_/D vssd1 vssd1 vccd1 vccd1 _15695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14646_ _16430_/Q _14756_/B _14655_/C vssd1 vssd1 vccd1 vccd1 _14646_/X sky130_fd_sc_hd__and3_1
X_11858_ _11891_/C vssd1 vssd1 vccd1 vccd1 _11897_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_33_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10809_ _10809_/A _10809_/B _10814_/B vssd1 vssd1 vccd1 vccd1 _15882_/D sky130_fd_sc_hd__nor3_1
XANTENNA_19 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _11901_/A _11795_/C vssd1 vssd1 vccd1 vccd1 _11789_/X sky130_fd_sc_hd__or2_1
X_14577_ _14575_/Y _14576_/X _14571_/C _14572_/C vssd1 vssd1 vccd1 vccd1 _14579_/B
+ sky130_fd_sc_hd__o211ai_1
X_16316_ _16346_/CLK _16316_/D vssd1 vssd1 vccd1 vccd1 _16316_/Q sky130_fd_sc_hd__dfxtp_1
X_13528_ _14220_/A vssd1 vssd1 vccd1 vccd1 _14092_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16247_ _16261_/CLK _16247_/D vssd1 vssd1 vccd1 vccd1 _16247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13459_ _16257_/Q _13573_/B _13459_/C vssd1 vssd1 vccd1 vccd1 _13459_/Y sky130_fd_sc_hd__nand3_1
X_16178_ _16237_/CLK _16178_/D vssd1 vssd1 vccd1 vccd1 _16178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15129_ _16508_/Q _15129_/B _15135_/C vssd1 vssd1 vccd1 vccd1 _15131_/C sky130_fd_sc_hd__nand3_1
XFILLER_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07951_ _15876_/Q vssd1 vssd1 vccd1 vccd1 _10675_/C sky130_fd_sc_hd__clkinv_2
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07882_ _07882_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _08132_/A sky130_fd_sc_hd__nand2_4
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09621_ _09953_/A vssd1 vssd1 vccd1 vccd1 _09718_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09552_ _09546_/C _09547_/C _09549_/Y _09556_/A vssd1 vssd1 vccd1 vccd1 _09556_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_83_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08503_ _08540_/B _08503_/B vssd1 vssd1 vccd1 vccd1 _08537_/A sky130_fd_sc_hd__and2_2
X_09483_ _09438_/X _09481_/B _09431_/X vssd1 vssd1 vccd1 vccd1 _09483_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08434_ _08344_/A _08344_/B _08433_/X vssd1 vssd1 vccd1 vccd1 _08476_/A sky130_fd_sc_hd__a21bo_1
XFILLER_51_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08365_ _08365_/A _08365_/B vssd1 vssd1 vccd1 vccd1 _08366_/B sky130_fd_sc_hd__xor2_2
XFILLER_149_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ _09987_/C _08296_/B vssd1 vssd1 vccd1 vccd1 _08296_/X sky130_fd_sc_hd__or2_1
XFILLER_3_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09819_ _09951_/A _09819_/B _09819_/C vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__and3_1
XFILLER_47_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _12823_/C _12824_/C _12826_/Y _12828_/X vssd1 vssd1 vccd1 vccd1 _12831_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_27_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _16159_/Q _12818_/B _12770_/C vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__and3_1
XFILLER_15_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14624_/A sky130_fd_sc_hd__buf_2
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11993_/A vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _16570_/CLK _15480_/D vssd1 vssd1 vccd1 vccd1 _15480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _16149_/Q _12798_/B _12692_/C vssd1 vssd1 vccd1 vccd1 _12701_/B sky130_fd_sc_hd__and3_1
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _16002_/Q _11648_/C _11591_/X vssd1 vssd1 vccd1 vccd1 _11643_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14484_/A _14431_/B _14435_/B vssd1 vssd1 vccd1 vccd1 _16395_/D sky130_fd_sc_hd__nor3_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11574_ _11594_/C vssd1 vssd1 vccd1 vccd1 _11607_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14362_ _14362_/A vssd1 vssd1 vccd1 vccd1 _16385_/D sky130_fd_sc_hd__clkbuf_1
X_16101_ _16554_/Q _16101_/D vssd1 vssd1 vccd1 vccd1 _16101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10525_ _10469_/X _10518_/B _10521_/B _10524_/Y vssd1 vssd1 vccd1 vccd1 _15829_/D
+ sky130_fd_sc_hd__o31a_1
X_13313_ _13313_/A _13313_/B vssd1 vssd1 vccd1 vccd1 _13314_/B sky130_fd_sc_hd__nor2_1
X_14293_ _14293_/A vssd1 vssd1 vccd1 vccd1 _16375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16032_ _16118_/CLK _16032_/D vssd1 vssd1 vccd1 vccd1 _16032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13244_ _13240_/Y _13241_/X _13243_/Y _13238_/C vssd1 vssd1 vccd1 vccd1 _13246_/B
+ sky130_fd_sc_hd__o211ai_1
X_10456_ _10456_/A vssd1 vssd1 vccd1 vccd1 _10652_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13175_ _13175_/A vssd1 vssd1 vccd1 vccd1 _16216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10387_ _15809_/Q _10388_/C _10243_/X vssd1 vssd1 vccd1 vccd1 _10387_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _12126_/A _12135_/B vssd1 vssd1 vccd1 vccd1 _12128_/A sky130_fd_sc_hd__or2_1
XFILLER_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12057_ _12057_/A vssd1 vssd1 vccd1 vccd1 _16058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11008_ _15911_/Q _11045_/C _10951_/X vssd1 vssd1 vccd1 vccd1 _11010_/B sky130_fd_sc_hd__a21oi_1
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15816_ _16595_/CLK _15816_/D vssd1 vssd1 vccd1 vccd1 _15816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15747_ _15812_/CLK _15747_/D vssd1 vssd1 vccd1 vccd1 _15747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12959_ _13242_/A vssd1 vssd1 vccd1 vccd1 _13187_/B sky130_fd_sc_hd__buf_2
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ _15791_/CLK _15678_/D vssd1 vssd1 vccd1 vccd1 _15678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14629_ _14629_/A _14629_/B _14629_/C vssd1 vssd1 vccd1 vccd1 _14630_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08150_ _10076_/C _08022_/B _08149_/X vssd1 vssd1 vccd1 vccd1 _08195_/A sky130_fd_sc_hd__o21ai_1
XFILLER_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ _15525_/Q _15507_/Q vssd1 vssd1 vccd1 vccd1 _08082_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _15532_/Q _08991_/C _08859_/X vssd1 vssd1 vccd1 vccd1 _08983_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ _16574_/Q vssd1 vssd1 vccd1 vccd1 _11798_/A sky130_fd_sc_hd__clkinv_4
XFILLER_29_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ _15732_/Q vssd1 vssd1 vccd1 vccd1 _09905_/C sky130_fd_sc_hd__clkinv_2
XFILLER_113_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _09604_/A vssd1 vssd1 vccd1 vccd1 _09604_/X sky130_fd_sc_hd__buf_2
X_07796_ _07799_/A vssd1 vssd1 vccd1 vccd1 _07796_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09535_ _09535_/A _09535_/B vssd1 vssd1 vccd1 vccd1 _15641_/D sky130_fd_sc_hd__nor2_1
X_09466_ _15631_/Q _09641_/B _09472_/C vssd1 vssd1 vccd1 vccd1 _09468_/B sky130_fd_sc_hd__and3_1
X_08417_ _15291_/A _08418_/B vssd1 vssd1 vccd1 vccd1 _08419_/A sky130_fd_sc_hd__or2_1
X_09397_ _09396_/X _10526_/A _09390_/B _08554_/A vssd1 vssd1 vccd1 vccd1 _09398_/B
+ sky130_fd_sc_hd__a31o_1
X_08348_ _08348_/A _08227_/A vssd1 vssd1 vccd1 vccd1 _08348_/X sky130_fd_sc_hd__or2b_1
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08279_ _08279_/A _08279_/B vssd1 vssd1 vccd1 vccd1 _08400_/A sky130_fd_sc_hd__xnor2_4
XFILLER_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10310_ _10308_/Y _10304_/C _10306_/Y _10315_/A vssd1 vssd1 vccd1 vccd1 _10315_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11290_ _11322_/C vssd1 vssd1 vccd1 vccd1 _11328_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10241_ _10250_/A _10241_/B _10241_/C vssd1 vssd1 vccd1 vccd1 _10242_/A sky130_fd_sc_hd__and3_1
XFILLER_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10172_ _10178_/C vssd1 vssd1 vccd1 vccd1 _10190_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14980_ _16483_/Q _14982_/C _14979_/X vssd1 vssd1 vccd1 vccd1 _14980_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_120_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13931_ _13931_/A _13931_/B vssd1 vssd1 vccd1 vccd1 _13933_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16643__48 vssd1 vssd1 vccd1 vccd1 _16643__48/HI _16719_/A sky130_fd_sc_hd__conb_1
X_13862_ _16315_/Q _13914_/B _13869_/C vssd1 vssd1 vccd1 vccd1 _13862_/X sky130_fd_sc_hd__and3_1
XFILLER_47_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15601_ _16551_/CLK _15601_/D vssd1 vssd1 vccd1 vccd1 _15601_/Q sky130_fd_sc_hd__dfxtp_1
X_12813_ _16592_/Q vssd1 vssd1 vccd1 vccd1 _12828_/C sky130_fd_sc_hd__inv_2
X_16581_ _16595_/CLK _16581_/D vssd1 vssd1 vccd1 vccd1 _16581_/Q sky130_fd_sc_hd__dfxtp_1
X_13793_ _16305_/Q _13900_/B _13793_/C vssd1 vssd1 vccd1 vccd1 _13793_/X sky130_fd_sc_hd__and3_1
XFILLER_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15532_ _16551_/CLK _15532_/D vssd1 vssd1 vccd1 vccd1 _15532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _16157_/Q _12745_/C _12575_/X vssd1 vssd1 vccd1 vccd1 _12746_/A sky130_fd_sc_hd__a21oi_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15463_ _16551_/CLK _15463_/D vssd1 vssd1 vccd1 vccd1 _15463_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _16147_/Q _12685_/C _12619_/X vssd1 vssd1 vccd1 vccd1 _12675_/Y sky130_fd_sc_hd__a21oi_1
X_14414_ _16393_/Q _14414_/B _14414_/C vssd1 vssd1 vccd1 vccd1 _14414_/Y sky130_fd_sc_hd__nand3_1
X_11626_ _11648_/C vssd1 vssd1 vccd1 vccd1 _11662_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15394_ _16053_/Q _16052_/Q _16051_/Q _15391_/X vssd1 vssd1 vccd1 vccd1 _16577_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14345_ _16384_/Q _14569_/B _14351_/C vssd1 vssd1 vccd1 vccd1 _14347_/C sky130_fd_sc_hd__nand3_1
XFILLER_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11557_ _11555_/Y _11547_/C _11550_/Y _11562_/A vssd1 vssd1 vccd1 vccd1 _11562_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10508_ _15829_/Q _10517_/C _10454_/X vssd1 vssd1 vccd1 vccd1 _10508_/Y sky130_fd_sc_hd__a21oi_1
X_11488_ _15978_/Q _11488_/B _11494_/C vssd1 vssd1 vccd1 vccd1 _11488_/Y sky130_fd_sc_hd__nand3_1
X_14276_ _14276_/A _14276_/B _14276_/C vssd1 vssd1 vccd1 vccd1 _14277_/C sky130_fd_sc_hd__or3_1
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _16118_/CLK _16015_/D vssd1 vssd1 vccd1 vccd1 _16015_/Q sky130_fd_sc_hd__dfxtp_1
X_13227_ _16225_/Q _13235_/C _13169_/X vssd1 vssd1 vccd1 vccd1 _13227_/Y sky130_fd_sc_hd__a21oi_1
X_10439_ _15818_/Q _10440_/C _10243_/X vssd1 vssd1 vccd1 vccd1 _10439_/Y sky130_fd_sc_hd__a21oi_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _16215_/Q _13199_/C _12933_/X vssd1 vssd1 vccd1 vccd1 _13161_/B sky130_fd_sc_hd__a21oi_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12109_ _13242_/A vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__clkbuf_2
X_13089_ _13087_/A _13087_/B _13088_/X vssd1 vssd1 vccd1 vccd1 _16204_/D sky130_fd_sc_hd__a21oi_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09320_ _15601_/Q _09448_/B _09320_/C vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__and3_1
X_09251_ _09267_/C vssd1 vssd1 vccd1 vccd1 _09286_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_08202_ _11964_/A _07983_/B _07982_/B vssd1 vssd1 vccd1 vccd1 _08204_/C sky130_fd_sc_hd__o21a_1
X_09182_ _09182_/A vssd1 vssd1 vccd1 vccd1 _15572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08133_ _13097_/A _07889_/B _08132_/X vssd1 vssd1 vccd1 vccd1 _08333_/B sky130_fd_sc_hd__o21a_1
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08064_ _08064_/A _08064_/B vssd1 vssd1 vccd1 vccd1 _08065_/B sky130_fd_sc_hd__nand2_2
XFILLER_134_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08966_ _08796_/X _08965_/A _08927_/X vssd1 vssd1 vccd1 vccd1 _08966_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07917_ _07917_/A _07917_/B vssd1 vssd1 vccd1 vccd1 _07949_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08897_ _08898_/B _08898_/C _08898_/A vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07848_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07848_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07779_ _07780_/A vssd1 vssd1 vccd1 vccd1 _07779_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09518_ _15262_/B vssd1 vssd1 vccd1 vccd1 _09692_/B sky130_fd_sc_hd__clkbuf_2
X_10790_ _11360_/A vssd1 vssd1 vccd1 vccd1 _11026_/B sky130_fd_sc_hd__buf_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09497_/A _09449_/B _09453_/A vssd1 vssd1 vccd1 vccd1 _15625_/D sky130_fd_sc_hd__nor3_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12460_ _12514_/A _12460_/B _12464_/B vssd1 vssd1 vccd1 vccd1 _16115_/D sky130_fd_sc_hd__nor3_1
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11411_ _11978_/A vssd1 vssd1 vccd1 vccd1 _11638_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_137_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12391_ _12391_/A vssd1 vssd1 vccd1 vccd1 _16105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11342_ _11375_/C vssd1 vssd1 vccd1 vccd1 _11381_/C sky130_fd_sc_hd__clkbuf_2
X_14130_ _14145_/A _14130_/B _14130_/C vssd1 vssd1 vccd1 vccd1 _14131_/A sky130_fd_sc_hd__and3_1
XFILLER_138_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11273_ _11379_/A _11273_/B _11277_/B vssd1 vssd1 vccd1 vccd1 _15947_/D sky130_fd_sc_hd__nor3_1
X_14061_ _16343_/Q _14101_/C _14060_/X vssd1 vssd1 vccd1 vccd1 _14063_/B sky130_fd_sc_hd__a21oi_1
XFILLER_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10224_ _10716_/A vssd1 vssd1 vccd1 vccd1 _10224_/X sky130_fd_sc_hd__clkbuf_2
X_13012_ _13019_/A _13012_/B _13012_/C vssd1 vssd1 vccd1 vccd1 _13013_/A sky130_fd_sc_hd__and3_1
XFILLER_133_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10155_ _10153_/Y _10145_/C _10147_/Y _10160_/A vssd1 vssd1 vccd1 vccd1 _10160_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10086_ _15755_/Q _10190_/B _10086_/C vssd1 vssd1 vccd1 vccd1 _10086_/X sky130_fd_sc_hd__and3_1
X_14963_ _14995_/C vssd1 vssd1 vccd1 vccd1 _15001_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16702_ _16702_/A _07802_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13914_ _16323_/Q _13914_/B _13923_/C vssd1 vssd1 vccd1 vccd1 _13914_/X sky130_fd_sc_hd__and3_1
XFILLER_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14894_ _14896_/B _14896_/C _14669_/X vssd1 vssd1 vccd1 vccd1 _14897_/B sky130_fd_sc_hd__o21ai_1
XFILLER_35_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13845_ _13866_/A _13845_/B _13845_/C vssd1 vssd1 vccd1 vccd1 _13846_/A sky130_fd_sc_hd__and3_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16564_ _16570_/CLK _16564_/D vssd1 vssd1 vccd1 vccd1 _16564_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13776_ _13776_/A vssd1 vssd1 vccd1 vccd1 _16301_/D sky130_fd_sc_hd__clkbuf_1
X_10988_ _10984_/Y _10994_/A _10987_/Y _10981_/C vssd1 vssd1 vccd1 vccd1 _10990_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15515_ _16551_/CLK _15515_/D vssd1 vssd1 vccd1 vccd1 _15515_/Q sky130_fd_sc_hd__dfxtp_1
X_12727_ _12724_/Y _12725_/X _12726_/Y _12721_/C vssd1 vssd1 vccd1 vccd1 _12729_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_31_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16495_ _16607_/CLK _16495_/D vssd1 vssd1 vccd1 vccd1 _16495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15446_ _16570_/CLK _15446_/D vssd1 vssd1 vccd1 vccd1 _15446_/Q sky130_fd_sc_hd__dfxtp_2
X_12658_ _12659_/B _12659_/C _12659_/A vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__a21o_1
X_11609_ _11606_/Y _11615_/A _11608_/Y _11604_/C vssd1 vssd1 vccd1 vccd1 _11611_/B
+ sky130_fd_sc_hd__o211a_1
X_15377_ _15949_/Q _15948_/Q _15947_/Q _15372_/X vssd1 vssd1 vccd1 vccd1 _16564_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_117_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12589_ _16588_/Q vssd1 vssd1 vccd1 vccd1 _12607_/C sky130_fd_sc_hd__inv_2
XFILLER_11_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14328_ _14326_/A _14326_/B _14327_/X vssd1 vssd1 vccd1 vccd1 _16380_/D sky130_fd_sc_hd__a21oi_1
XFILLER_117_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14259_ _16372_/Q _14268_/C _14258_/X vssd1 vssd1 vccd1 vccd1 _14259_/Y sky130_fd_sc_hd__a21oi_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _10789_/B vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__buf_4
XFILLER_98_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _10414_/A vssd1 vssd1 vccd1 vccd1 _08921_/B sky130_fd_sc_hd__clkbuf_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08682_ _08682_/A vssd1 vssd1 vccd1 vccd1 _15464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09303_ _15058_/A vssd1 vssd1 vccd1 vccd1 _09750_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_139_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09234_ _09234_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09235_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09165_ _15358_/A _15358_/B _09165_/C vssd1 vssd1 vccd1 vccd1 _09167_/A sky130_fd_sc_hd__and3_1
XFILLER_119_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08116_ _09448_/C _08116_/B vssd1 vssd1 vccd1 vccd1 _08116_/X sky130_fd_sc_hd__or2_1
XFILLER_147_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ _15557_/Q _15332_/B _09099_/C vssd1 vssd1 vccd1 vccd1 _09101_/A sky130_fd_sc_hd__and3_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08047_ _10029_/C _08047_/B vssd1 vssd1 vccd1 vccd1 _08048_/B sky130_fd_sc_hd__xnor2_4
XFILLER_116_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09998_ _15738_/Q _09998_/B _09998_/C vssd1 vssd1 vccd1 vccd1 _10004_/A sky130_fd_sc_hd__and3_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08949_ _08949_/A _08949_/B vssd1 vssd1 vccd1 vccd1 _08951_/A sky130_fd_sc_hd__or2_1
XFILLER_57_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11960_ _12018_/A _11960_/B _11960_/C vssd1 vssd1 vccd1 vccd1 _11961_/C sky130_fd_sc_hd__or3_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10911_ _10911_/A vssd1 vssd1 vccd1 vccd1 _15896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11891_ _16036_/Q _11891_/B _11891_/C vssd1 vssd1 vccd1 vccd1 _11899_/A sky130_fd_sc_hd__and3_1
XFILLER_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13630_ _16283_/Q _13639_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13630_/Y sky130_fd_sc_hd__a21oi_1
X_10842_ _12886_/A vssd1 vssd1 vccd1 vccd1 _11978_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13561_ _13561_/A _13561_/B _13561_/C vssd1 vssd1 vccd1 vccd1 _13562_/C sky130_fd_sc_hd__nand3_1
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10773_ _10809_/A _10773_/B _10777_/A vssd1 vssd1 vccd1 vccd1 _15877_/D sky130_fd_sc_hd__nor3_1
XFILLER_9_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15300_ _15300_/A vssd1 vssd1 vccd1 vccd1 _15301_/B sky130_fd_sc_hd__inv_2
X_12512_ _12507_/Y _12518_/A _12511_/Y _12505_/C vssd1 vssd1 vccd1 vccd1 _12514_/B
+ sky130_fd_sc_hd__o211a_1
X_16280_ _16533_/Q _16280_/D vssd1 vssd1 vccd1 vccd1 _16280_/Q sky130_fd_sc_hd__dfxtp_1
X_13492_ _13507_/C vssd1 vssd1 vccd1 vccd1 _13514_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15231_ _16525_/Q _15267_/C _08843_/A vssd1 vssd1 vccd1 vccd1 _15233_/B sky130_fd_sc_hd__a21oi_1
XFILLER_100_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12443_ _16113_/Q _12443_/B _12443_/C vssd1 vssd1 vccd1 vccd1 _12443_/Y sky130_fd_sc_hd__nand3_1
XFILLER_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15162_ _15162_/A _15169_/B vssd1 vssd1 vccd1 vccd1 _15164_/A sky130_fd_sc_hd__or2_1
X_12374_ _16104_/Q _12600_/B _12380_/C vssd1 vssd1 vccd1 vccd1 _12376_/C sky130_fd_sc_hd__nand3_1
X_14113_ _14113_/A vssd1 vssd1 vccd1 vccd1 _14127_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11325_ _11323_/Y _11319_/C _11321_/Y _11330_/A vssd1 vssd1 vccd1 vccd1 _11330_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15093_ _15100_/A _15093_/B _15093_/C vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__and3_1
XFILLER_125_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11256_ _11264_/A _11256_/B _11256_/C vssd1 vssd1 vccd1 vccd1 _11257_/A sky130_fd_sc_hd__and3_1
X_14044_ _16341_/Q _14207_/B _14044_/C vssd1 vssd1 vccd1 vccd1 _14053_/B sky130_fd_sc_hd__and3_1
XFILLER_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10207_ _10510_/A vssd1 vssd1 vccd1 vccd1 _10458_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_122_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11187_ _11187_/A vssd1 vssd1 vccd1 vccd1 _15935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10138_ _10393_/A vssd1 vssd1 vccd1 vccd1 _10138_/X sky130_fd_sc_hd__buf_2
X_15995_ _16005_/CLK _15995_/D vssd1 vssd1 vccd1 vccd1 _15995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10069_ _15704_/Q _15703_/Q _15702_/Q _09982_/X vssd1 vssd1 vccd1 vccd1 _15750_/D
+ sky130_fd_sc_hd__o31a_1
X_14946_ _16477_/Q _14947_/C _14828_/X vssd1 vssd1 vccd1 vccd1 _14948_/A sky130_fd_sc_hd__a21oi_1
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14877_ _14875_/Y _14870_/C _14873_/Y _14874_/X vssd1 vssd1 vccd1 vccd1 _14878_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16616_ input11/X _16616_/D vssd1 vssd1 vccd1 vccd1 _16616_/Q sky130_fd_sc_hd__dfxtp_1
X_13828_ _13881_/A vssd1 vssd1 vccd1 vccd1 _13866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16547_ _16551_/CLK _16547_/D vssd1 vssd1 vccd1 vccd1 _16547_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ _16300_/Q _13869_/B _13759_/C vssd1 vssd1 vccd1 vccd1 _13767_/A sky130_fd_sc_hd__and3_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16478_ _16607_/CLK _16478_/D vssd1 vssd1 vccd1 vccd1 _16478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15429_ _16277_/Q _16276_/Q _16275_/Q _15428_/X vssd1 vssd1 vccd1 vccd1 _16605_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_117_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09921_ _09921_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _09921_/X sky130_fd_sc_hd__or2_1
X_16679__84 vssd1 vssd1 vccd1 vccd1 _16679__84/HI _16755_/A sky130_fd_sc_hd__conb_1
XFILLER_125_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09852_ _09846_/B _09849_/B _09125_/A vssd1 vssd1 vccd1 vccd1 _09853_/B sky130_fd_sc_hd__o21a_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08803_ _15494_/Q _08845_/B _08807_/C vssd1 vssd1 vccd1 vccd1 _08809_/A sky130_fd_sc_hd__and3_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09783_ _09781_/X _09783_/B vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__and2b_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08734_ _08734_/A _08734_/B vssd1 vssd1 vccd1 vccd1 _08735_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _08661_/X _08656_/A _08664_/Y vssd1 vssd1 vccd1 vccd1 _15461_/D sky130_fd_sc_hd__o21a_1
XFILLER_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _13085_/A vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__buf_4
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09217_ _10900_/B vssd1 vssd1 vccd1 vccd1 _09629_/A sky130_fd_sc_hd__buf_4
XFILLER_148_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09148_ _09148_/A _09148_/B _09152_/B vssd1 vssd1 vccd1 vccd1 _15564_/D sky130_fd_sc_hd__nor3_1
XFILLER_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09079_ _09076_/X _09071_/B _09074_/B _09078_/Y vssd1 vssd1 vccd1 vccd1 _15548_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11110_ _11148_/A _11110_/B _11110_/C vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__and3_1
XFILLER_123_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12090_ _12113_/A _12090_/B _12090_/C vssd1 vssd1 vccd1 vccd1 _12091_/A sky130_fd_sc_hd__and3_1
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11041_ _11038_/Y _11047_/A _11040_/Y _11036_/C vssd1 vssd1 vccd1 vccd1 _11043_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14800_ _16455_/Q _15027_/B _14800_/C vssd1 vssd1 vccd1 vccd1 _14800_/X sky130_fd_sc_hd__and3_1
X_15780_ _16595_/CLK _15780_/D vssd1 vssd1 vccd1 vccd1 _15780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12992_ _16191_/Q _13102_/B _13001_/C vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__and3_1
XFILLER_18_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14731_ _14764_/C vssd1 vssd1 vccd1 vccd1 _14770_/C sky130_fd_sc_hd__clkbuf_2
X_11943_ _12225_/A vssd1 vssd1 vccd1 vccd1 _12173_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14662_ _16432_/Q _14770_/B _14662_/C vssd1 vssd1 vccd1 vccd1 _14671_/B sky130_fd_sc_hd__and3_1
X_11874_ _13288_/A vssd1 vssd1 vccd1 vccd1 _13006_/A sky130_fd_sc_hd__buf_4
X_16401_ input11/X _16401_/D vssd1 vssd1 vccd1 vccd1 _16401_/Q sky130_fd_sc_hd__dfxtp_1
X_13613_ _13613_/A _13613_/B _13613_/C vssd1 vssd1 vccd1 vccd1 _13614_/C sky130_fd_sc_hd__nand3_1
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10825_ _10825_/A vssd1 vssd1 vccd1 vccd1 _15884_/D sky130_fd_sc_hd__clkbuf_1
X_14593_ _14591_/Y _14586_/C _14589_/Y _14590_/X vssd1 vssd1 vccd1 vccd1 _14594_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16332_ _16346_/CLK _16332_/D vssd1 vssd1 vccd1 vccd1 _16332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13544_ _13598_/A vssd1 vssd1 vccd1 vccd1 _13583_/A sky130_fd_sc_hd__clkbuf_2
X_10756_ _10756_/A _10756_/B vssd1 vssd1 vccd1 vccd1 _10758_/A sky130_fd_sc_hd__or2_1
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16263_ _16533_/Q _16263_/D vssd1 vssd1 vccd1 vccd1 _16263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13475_ _13472_/Y _13481_/A _13474_/Y _13470_/C vssd1 vssd1 vccd1 vccd1 _13477_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10687_ _10681_/C _10682_/C _10684_/Y _10685_/X vssd1 vssd1 vccd1 vccd1 _10688_/C
+ sky130_fd_sc_hd__a211o_1
X_15214_ _16522_/Q _15215_/C _10812_/B vssd1 vssd1 vccd1 vccd1 _15216_/A sky130_fd_sc_hd__a21oi_1
X_12426_ _16111_/Q _12535_/B _12435_/C vssd1 vssd1 vccd1 vccd1 _12431_/A sky130_fd_sc_hd__and3_1
X_16194_ _16555_/Q _16194_/D vssd1 vssd1 vccd1 vccd1 _16194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15145_ _15152_/A _15145_/B _15145_/C vssd1 vssd1 vccd1 vccd1 _15146_/A sky130_fd_sc_hd__and3_1
XFILLER_126_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12357_ _12355_/A _12355_/B _12356_/X vssd1 vssd1 vccd1 vccd1 _16100_/D sky130_fd_sc_hd__a21oi_1
XFILLER_5_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11308_ _15954_/Q _11359_/B _11309_/C vssd1 vssd1 vccd1 vccd1 _11308_/X sky130_fd_sc_hd__and3_1
X_15076_ _16499_/Q _15083_/C _14851_/X vssd1 vssd1 vccd1 vccd1 _15079_/B sky130_fd_sc_hd__a21o_1
XFILLER_114_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12288_ _16091_/Q _12347_/B _12296_/C vssd1 vssd1 vccd1 vccd1 _12288_/Y sky130_fd_sc_hd__nand3_1
X_14027_ _14035_/A _14027_/B _14027_/C vssd1 vssd1 vccd1 vccd1 _14028_/A sky130_fd_sc_hd__and3_1
X_11239_ _12373_/A vssd1 vssd1 vccd1 vccd1 _11465_/B sky130_fd_sc_hd__buf_2
XFILLER_68_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15978_ _16005_/CLK _15978_/D vssd1 vssd1 vccd1 vccd1 _15978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14929_ _14929_/A vssd1 vssd1 vccd1 vccd1 _16473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08450_ _08355_/A _08355_/B _08359_/B vssd1 vssd1 vccd1 vccd1 _08450_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ _08241_/A _08241_/B _08380_/Y vssd1 vssd1 vccd1 vccd1 _08384_/A sky130_fd_sc_hd__o21ai_4
XFILLER_51_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09002_ _09002_/A _09002_/B vssd1 vssd1 vccd1 vccd1 _15531_/D sky130_fd_sc_hd__nor2_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09904_ _15718_/Q _09925_/C _09714_/X vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__a21oi_1
XFILLER_58_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09835_ _15703_/Q _09845_/C _10009_/B vssd1 vssd1 vccd1 vccd1 _09835_/Y sky130_fd_sc_hd__a21oi_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _09766_/A _09766_/B _09766_/C vssd1 vssd1 vccd1 vccd1 _09767_/C sky130_fd_sc_hd__nand3_1
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08717_ _15476_/Q _08732_/C _08576_/X vssd1 vssd1 vccd1 vccd1 _08719_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _09691_/Y _09692_/X _09694_/B vssd1 vssd1 vccd1 vccd1 _09700_/B sky130_fd_sc_hd__o21a_1
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _12574_/A vssd1 vssd1 vccd1 vccd1 _14828_/A sky130_fd_sc_hd__buf_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _15367_/B _08579_/B _08592_/A vssd1 vssd1 vccd1 vccd1 _15454_/D sky130_fd_sc_hd__nor3_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10676_/A _10610_/B _10614_/B vssd1 vssd1 vccd1 vccd1 _15845_/D sky130_fd_sc_hd__nor3_1
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11590_ _11590_/A vssd1 vssd1 vccd1 vccd1 _15992_/D sky130_fd_sc_hd__clkbuf_1
X_10541_ _10541_/A _10541_/B _10541_/C vssd1 vssd1 vccd1 vccd1 _10542_/C sky130_fd_sc_hd__nand3_1
XFILLER_128_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _13260_/A _13260_/B vssd1 vssd1 vccd1 vccd1 _13266_/C sky130_fd_sc_hd__nor2_1
XFILLER_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10472_ _10469_/X _10464_/B _10467_/B _10471_/Y vssd1 vssd1 vccd1 vccd1 _15820_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12211_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12443_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_136_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13191_ _13191_/A vssd1 vssd1 vccd1 vccd1 _16218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12142_ _16071_/Q _12179_/C _12081_/X vssd1 vssd1 vccd1 vccd1 _12144_/B sky130_fd_sc_hd__a21oi_1
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12073_ _12924_/A vssd1 vssd1 vccd1 vccd1 _12304_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15901_ _16553_/Q _15901_/D vssd1 vssd1 vccd1 vccd1 _15901_/Q sky130_fd_sc_hd__dfxtp_1
X_11024_ _15914_/Q _11026_/C _11023_/X vssd1 vssd1 vccd1 vccd1 _11024_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832_ _16595_/CLK _15832_/D vssd1 vssd1 vccd1 vccd1 _15832_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15763_ _15791_/CLK _15763_/D vssd1 vssd1 vccd1 vccd1 _15763_/Q sky130_fd_sc_hd__dfxtp_1
X_12975_ _16189_/Q _13082_/B _12975_/C vssd1 vssd1 vccd1 vccd1 _12984_/B sky130_fd_sc_hd__and3_1
XFILLER_18_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14714_ _14768_/A _14714_/B _14718_/B vssd1 vssd1 vccd1 vccd1 _16439_/D sky130_fd_sc_hd__nor3_1
X_11926_ _11926_/A vssd1 vssd1 vccd1 vccd1 _16040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15694_ _15791_/CLK _15694_/D vssd1 vssd1 vccd1 vccd1 _15694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14645_ _16430_/Q _14655_/C _14588_/X vssd1 vssd1 vccd1 vccd1 _14645_/Y sky130_fd_sc_hd__a21oi_1
X_11857_ _11878_/C vssd1 vssd1 vccd1 vccd1 _11891_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10808_ _10806_/Y _10801_/C _10803_/Y _10814_/A vssd1 vssd1 vccd1 vccd1 _10814_/B
+ sky130_fd_sc_hd__a211oi_1
X_14576_ _16419_/Q _14742_/B _14576_/C vssd1 vssd1 vccd1 vccd1 _14576_/X sky130_fd_sc_hd__and3_1
X_11788_ _11788_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11795_/C sky130_fd_sc_hd__nor2_1
X_16315_ _16346_/CLK _16315_/D vssd1 vssd1 vccd1 vccd1 _16315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13527_ _13527_/A vssd1 vssd1 vccd1 vccd1 _16266_/D sky130_fd_sc_hd__clkbuf_1
X_10739_ _10739_/A vssd1 vssd1 vccd1 vccd1 _15870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16246_ _16261_/CLK _16246_/D vssd1 vssd1 vccd1 vccd1 _16246_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13458_ _16258_/Q _13623_/B _13459_/C vssd1 vssd1 vccd1 vccd1 _13458_/X sky130_fd_sc_hd__and3_1
X_12409_ _16109_/Q _12516_/B _12409_/C vssd1 vssd1 vccd1 vccd1 _12418_/B sky130_fd_sc_hd__and3_1
X_16177_ _16237_/CLK _16177_/D vssd1 vssd1 vccd1 vccd1 _16177_/Q sky130_fd_sc_hd__dfxtp_1
X_13389_ _13412_/A _13389_/B _13389_/C vssd1 vssd1 vccd1 vccd1 _13390_/A sky130_fd_sc_hd__and3_1
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15128_ _16508_/Q _15135_/C _10956_/A vssd1 vssd1 vccd1 vccd1 _15131_/B sky130_fd_sc_hd__a21o_1
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16649__54 vssd1 vssd1 vccd1 vccd1 _16649__54/HI _16725_/A sky130_fd_sc_hd__conb_1
X_07950_ _15750_/Q vssd1 vssd1 vccd1 vccd1 _09802_/C sky130_fd_sc_hd__clkinv_4
X_15059_ _15059_/A _15059_/B vssd1 vssd1 vccd1 vccd1 _15064_/C sky130_fd_sc_hd__nor2_1
XFILLER_102_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07881_ _16442_/Q _07881_/B _08129_/A vssd1 vssd1 vccd1 vccd1 _08129_/B sky130_fd_sc_hd__nand3_2
XFILLER_96_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ _15650_/Q _15649_/Q _15648_/Q _09536_/X vssd1 vssd1 vccd1 vccd1 _15660_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_96_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09551_ _09549_/Y _09556_/A _09546_/C _09547_/C vssd1 vssd1 vccd1 vccd1 _09553_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08502_ _08502_/A _08502_/B _08502_/C vssd1 vssd1 vccd1 vccd1 _08503_/B sky130_fd_sc_hd__nand3_1
X_09482_ _09291_/X _09480_/B _09481_/Y vssd1 vssd1 vccd1 vccd1 _15630_/D sky130_fd_sc_hd__o21a_1
XFILLER_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08433_ _08433_/A _08345_/A vssd1 vssd1 vccd1 vccd1 _08433_/X sky130_fd_sc_hd__or2b_1
XFILLER_51_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08364_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _08365_/B sky130_fd_sc_hd__nor2_1
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08295_ _08295_/A vssd1 vssd1 vccd1 vccd1 _09178_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09818_ _09809_/C _09810_/C _09814_/Y _09816_/X vssd1 vssd1 vccd1 vccd1 _09819_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09749_ _09749_/A vssd1 vssd1 vccd1 vccd1 _09749_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _16159_/Q _12798_/C _12650_/X vssd1 vssd1 vccd1 vccd1 _12762_/B sky130_fd_sc_hd__a21oi_1
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _16011_/Q _11721_/C _11485_/X vssd1 vssd1 vccd1 vccd1 _11711_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12691_ _16149_/Q _12692_/C _12575_/X vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__a21oi_1
XFILLER_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14428_/Y _14424_/C _14426_/Y _14435_/A vssd1 vssd1 vccd1 vccd1 _14435_/B
+ sky130_fd_sc_hd__a211oi_1
X_11642_ _11642_/A vssd1 vssd1 vccd1 vccd1 _16000_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _14369_/A _14361_/B _14361_/C vssd1 vssd1 vccd1 vccd1 _14362_/A sky130_fd_sc_hd__and3_1
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11573_ _11586_/C vssd1 vssd1 vccd1 vccd1 _11594_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_128_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16100_ _16554_/Q _16100_/D vssd1 vssd1 vccd1 vccd1 _16100_/Q sky130_fd_sc_hd__dfxtp_1
X_13312_ _13312_/A _13319_/B vssd1 vssd1 vccd1 vccd1 _13314_/A sky130_fd_sc_hd__or2_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10524_ _10573_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10524_/Y sky130_fd_sc_hd__nor2_1
X_14292_ _14314_/A _14292_/B _14292_/C vssd1 vssd1 vccd1 vccd1 _14293_/A sky130_fd_sc_hd__and3_1
X_16031_ _16118_/CLK _16031_/D vssd1 vssd1 vccd1 vccd1 _16031_/Q sky130_fd_sc_hd__dfxtp_1
X_13243_ _16226_/Q _13467_/B _13250_/C vssd1 vssd1 vccd1 vccd1 _13243_/Y sky130_fd_sc_hd__nand3_1
X_10455_ _15820_/Q _10463_/C _10454_/X vssd1 vssd1 vccd1 vccd1 _10455_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13174_ _13190_/A _13174_/B _13174_/C vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__and3_1
X_10386_ _10386_/A vssd1 vssd1 vccd1 vccd1 _15806_/D sky130_fd_sc_hd__clkbuf_1
X_12125_ _16069_/Q _12232_/B _12125_/C vssd1 vssd1 vccd1 vccd1 _12135_/B sky130_fd_sc_hd__and3_1
XFILLER_69_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _12056_/A _12056_/B _12056_/C vssd1 vssd1 vccd1 vccd1 _12057_/A sky130_fd_sc_hd__and3_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _11039_/C vssd1 vssd1 vccd1 vccd1 _11045_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15815_ _16595_/CLK _15815_/D vssd1 vssd1 vccd1 vccd1 _15815_/Q sky130_fd_sc_hd__dfxtp_2
X_15746_ _15791_/CLK _15746_/D vssd1 vssd1 vccd1 vccd1 _15746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12958_ _16187_/Q _13068_/B _12967_/C vssd1 vssd1 vccd1 vccd1 _12958_/X sky130_fd_sc_hd__and3_1
X_11909_ _11922_/C vssd1 vssd1 vccd1 vccd1 _11930_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15677_ _15791_/CLK _15677_/D vssd1 vssd1 vccd1 vccd1 _15677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _16177_/Q _13053_/B _12889_/C vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__and3_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14628_ _14629_/B _14629_/C _14629_/A vssd1 vssd1 vccd1 vccd1 _14630_/B sky130_fd_sc_hd__a21o_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14559_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14576_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _15525_/Q _15507_/Q vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__or2_1
XFILLER_146_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16229_ _16237_/CLK _16229_/D vssd1 vssd1 vccd1 vccd1 _16229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08982_ _08982_/A vssd1 vssd1 vccd1 vccd1 _15527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07933_ _07933_/A _07933_/B vssd1 vssd1 vccd1 vccd1 _07945_/A sky130_fd_sc_hd__nor2_2
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07864_ _15714_/Q vssd1 vssd1 vccd1 vccd1 _09255_/C sky130_fd_sc_hd__inv_2
XFILLER_110_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09603_ _15659_/Q _09692_/B _09603_/C vssd1 vssd1 vccd1 vccd1 _09603_/X sky130_fd_sc_hd__and3_1
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07795_ _07799_/A vssd1 vssd1 vccd1 vccd1 _07795_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09534_ _09396_/X _09486_/X _09527_/B _09487_/X vssd1 vssd1 vccd1 vccd1 _09535_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09465_ _15255_/B vssd1 vssd1 vccd1 vccd1 _09641_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08416_ _15449_/Q _08490_/A vssd1 vssd1 vccd1 vccd1 _08418_/B sky130_fd_sc_hd__and2_1
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09396_ _09898_/A vssd1 vssd1 vccd1 vccd1 _09396_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08347_ _08194_/A _08194_/B _08346_/Y vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__a21o_2
XFILLER_149_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08278_ _08396_/A _08396_/B vssd1 vssd1 vccd1 vccd1 _08279_/B sky130_fd_sc_hd__xor2_4
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10240_ _10240_/A _10240_/B _10240_/C vssd1 vssd1 vccd1 vccd1 _10241_/C sky130_fd_sc_hd__nand3_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10171_ _15758_/Q _15757_/Q _15756_/Q _09982_/X vssd1 vssd1 vccd1 vccd1 _15768_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_79_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13930_ _13930_/A _13939_/B vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__or2_1
XFILLER_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13861_ _16315_/Q _13869_/C _13750_/X vssd1 vssd1 vccd1 vccd1 _13861_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15600_ _16570_/CLK _15600_/D vssd1 vssd1 vccd1 vccd1 _15600_/Q sky130_fd_sc_hd__dfxtp_2
X_12812_ _13377_/A vssd1 vssd1 vccd1 vccd1 _12936_/A sky130_fd_sc_hd__buf_2
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16580_ _16595_/CLK _16580_/D vssd1 vssd1 vccd1 vccd1 _16580_/Q sky130_fd_sc_hd__dfxtp_1
X_13792_ _16305_/Q _13800_/C _13736_/X vssd1 vssd1 vccd1 vccd1 _13792_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15531_ _16551_/CLK _15531_/D vssd1 vssd1 vccd1 vccd1 _15531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12796_/A _12743_/B _12747_/B vssd1 vssd1 vccd1 vccd1 _16155_/D sky130_fd_sc_hd__nor3_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15462_ _16551_/CLK _15462_/D vssd1 vssd1 vccd1 vccd1 _15462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12674_ _12674_/A vssd1 vssd1 vccd1 vccd1 _16145_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _16394_/Q _14464_/B _14414_/C vssd1 vssd1 vccd1 vccd1 _14413_/X sky130_fd_sc_hd__and3_1
X_11625_ _11638_/C vssd1 vssd1 vccd1 vccd1 _11648_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15393_ _16045_/Q _16044_/Q _16043_/Q _15391_/X vssd1 vssd1 vccd1 vccd1 _16576_/D
+ sky130_fd_sc_hd__o31a_1
X_14344_ _14911_/A vssd1 vssd1 vccd1 vccd1 _14569_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_129_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11556_ _11550_/Y _11562_/A _11555_/Y _11547_/C vssd1 vssd1 vccd1 vccd1 _11558_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10507_ _10507_/A vssd1 vssd1 vccd1 vccd1 _15826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14275_ _14276_/B _14276_/C _14108_/X vssd1 vssd1 vccd1 vccd1 _14277_/B sky130_fd_sc_hd__o21ai_1
X_11487_ _15979_/Q _11654_/B _11494_/C vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__and3_1
X_16014_ _16554_/Q _16014_/D vssd1 vssd1 vccd1 vccd1 _16014_/Q sky130_fd_sc_hd__dfxtp_2
X_13226_ _13226_/A vssd1 vssd1 vccd1 vccd1 _16223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10438_ _10438_/A vssd1 vssd1 vccd1 vccd1 _15815_/D sky130_fd_sc_hd__clkbuf_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13157_ _13193_/C vssd1 vssd1 vccd1 vccd1 _13199_/C sky130_fd_sc_hd__clkbuf_2
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _10363_/B _10366_/B _10164_/X vssd1 vssd1 vccd1 vccd1 _10370_/B sky130_fd_sc_hd__o21a_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12108_ _15247_/B vssd1 vssd1 vccd1 vccd1 _13242_/A sky130_fd_sc_hd__buf_4
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _13315_/A _13093_/C vssd1 vssd1 vccd1 vccd1 _13088_/X sky130_fd_sc_hd__or2_1
XFILLER_111_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12039_ _12037_/Y _12038_/X _12033_/C _12034_/C vssd1 vssd1 vccd1 vccd1 _12041_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15729_ _15812_/CLK _15729_/D vssd1 vssd1 vccd1 vccd1 _15729_/Q sky130_fd_sc_hd__dfxtp_1
X_09250_ _09255_/C vssd1 vssd1 vccd1 vccd1 _09267_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08201_ _11004_/A _08053_/B _08200_/X vssd1 vssd1 vccd1 vccd1 _08226_/A sky130_fd_sc_hd__o21ai_2
X_09181_ _09367_/A _09181_/B _09181_/C vssd1 vssd1 vccd1 vccd1 _09182_/A sky130_fd_sc_hd__and3_1
XFILLER_147_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08132_ _08132_/A _08132_/B vssd1 vssd1 vccd1 vccd1 _08132_/X sky130_fd_sc_hd__or2_1
XFILLER_147_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ _15633_/Q _15615_/Q vssd1 vssd1 vccd1 vccd1 _08064_/B sky130_fd_sc_hd__or2_1
XFILLER_134_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08965_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _15523_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07916_ _11572_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07917_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08896_ _15513_/Q _09016_/B _08896_/C vssd1 vssd1 vccd1 vccd1 _08898_/C sky130_fd_sc_hd__nand3_1
XFILLER_84_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07847_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07847_/Y sky130_fd_sc_hd__inv_2
X_07778_ _07780_/A vssd1 vssd1 vccd1 vccd1 _07778_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _09514_/A _09513_/Y _09514_/B vssd1 vssd1 vccd1 vccd1 _09517_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _15628_/Q _09448_/B _09448_/C vssd1 vssd1 vccd1 vccd1 _09453_/A sky130_fd_sc_hd__and3_1
XFILLER_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ _09378_/X _09377_/Y _10017_/A vssd1 vssd1 vccd1 vccd1 _09379_/Y sky130_fd_sc_hd__a21oi_1
X_11410_ _15969_/Q _11420_/C _11188_/X vssd1 vssd1 vccd1 vccd1 _11410_/Y sky130_fd_sc_hd__a21oi_1
X_12390_ _12398_/A _12390_/B _12390_/C vssd1 vssd1 vccd1 vccd1 _12391_/A sky130_fd_sc_hd__and3_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11341_ _11361_/C vssd1 vssd1 vccd1 vccd1 _11375_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14060_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14060_/X sky130_fd_sc_hd__clkbuf_2
X_11272_ _11270_/Y _11264_/C _11267_/Y _11277_/A vssd1 vssd1 vccd1 vccd1 _11277_/B
+ sky130_fd_sc_hd__a211oi_1
X_13011_ _13009_/Y _13004_/C _13007_/Y _13008_/X vssd1 vssd1 vccd1 vccd1 _13012_/C
+ sky130_fd_sc_hd__a211o_1
X_10223_ _10220_/X _10215_/B _10218_/B _10222_/Y vssd1 vssd1 vccd1 vccd1 _15775_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_121_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10154_ _10147_/Y _10160_/A _10153_/Y _10145_/C vssd1 vssd1 vccd1 vccd1 _10156_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14962_ _14982_/C vssd1 vssd1 vccd1 vccd1 _14995_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10085_ _15755_/Q _10086_/C _09813_/X vssd1 vssd1 vccd1 vccd1 _10085_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16701_ _16701_/A _07801_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
X_13913_ _16323_/Q _13923_/C _13750_/X vssd1 vssd1 vccd1 vccd1 _13913_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14893_ _15007_/A vssd1 vssd1 vccd1 vccd1 _14936_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13844_ _13844_/A _13844_/B _13844_/C vssd1 vssd1 vccd1 vccd1 _13845_/C sky130_fd_sc_hd__nand3_1
XFILLER_28_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16563_ _16570_/CLK _16563_/D vssd1 vssd1 vccd1 vccd1 _16563_/Q sky130_fd_sc_hd__dfxtp_2
X_13775_ _13811_/A _13775_/B _13775_/C vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__and3_1
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ _15907_/Q _11212_/B _10992_/C vssd1 vssd1 vccd1 vccd1 _10987_/Y sky130_fd_sc_hd__nand3_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12726_ _16153_/Q _12726_/B _12726_/C vssd1 vssd1 vccd1 vccd1 _12726_/Y sky130_fd_sc_hd__nand3_1
X_15514_ _16551_/CLK _15514_/D vssd1 vssd1 vccd1 vccd1 _15514_/Q sky130_fd_sc_hd__dfxtp_1
X_16494_ _16607_/CLK _16494_/D vssd1 vssd1 vccd1 vccd1 _16494_/Q sky130_fd_sc_hd__dfxtp_1
X_15445_ _16389_/Q _16388_/Q _16387_/Q _15440_/X vssd1 vssd1 vccd1 vccd1 _16619_/D
+ sky130_fd_sc_hd__o31a_1
X_12657_ _16144_/Q _12881_/B _12663_/C vssd1 vssd1 vccd1 vccd1 _12659_/C sky130_fd_sc_hd__nand3_1
XFILLER_129_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11608_ _15995_/Q _11780_/B _11613_/C vssd1 vssd1 vccd1 vccd1 _11608_/Y sky130_fd_sc_hd__nand3_1
X_15376_ _15941_/Q _15940_/Q _15939_/Q _15372_/X vssd1 vssd1 vccd1 vccd1 _16563_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12588_ _12588_/A vssd1 vssd1 vccd1 vccd1 _16133_/D sky130_fd_sc_hd__clkbuf_1
X_14327_ _14437_/A _14332_/C vssd1 vssd1 vccd1 vccd1 _14327_/X sky130_fd_sc_hd__or2_1
XFILLER_128_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11539_ _11547_/A _11539_/B _11539_/C vssd1 vssd1 vccd1 vccd1 _11540_/A sky130_fd_sc_hd__and3_1
XFILLER_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14258_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13209_ _13432_/A _13209_/B _13209_/C vssd1 vssd1 vccd1 vccd1 _13210_/C sky130_fd_sc_hd__or3_1
XFILLER_125_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14187_/Y _14182_/C _14184_/Y _14185_/X vssd1 vssd1 vccd1 vccd1 _14190_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _09164_/A vssd1 vssd1 vccd1 vccd1 _10414_/A sky130_fd_sc_hd__buf_4
XFILLER_100_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08681_ _15304_/A _08681_/B _08681_/C vssd1 vssd1 vccd1 vccd1 _08682_/A sky130_fd_sc_hd__and3_1
XFILLER_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09302_ input8/X vssd1 vssd1 vccd1 vccd1 _15058_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _09233_/A _09233_/B vssd1 vssd1 vccd1 vccd1 _09234_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09164_ _09164_/A vssd1 vssd1 vccd1 vccd1 _15358_/B sky130_fd_sc_hd__clkbuf_2
X_08115_ _09016_/C _08102_/B _08114_/Y vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__o21ai_4
X_09095_ _10285_/C vssd1 vssd1 vccd1 vccd1 _15332_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08046_ _08046_/A _08046_/B vssd1 vssd1 vccd1 vccd1 _08047_/B sky130_fd_sc_hd__nand2_2
XFILLER_150_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09997_ _15738_/Q _09998_/C _08604_/A vssd1 vssd1 vccd1 vccd1 _09997_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08948_ _15524_/Q _08991_/B _08948_/C vssd1 vssd1 vccd1 vccd1 _08949_/B sky130_fd_sc_hd__and3_1
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08879_ _08879_/A _08879_/B vssd1 vssd1 vccd1 vccd1 _15504_/D sky130_fd_sc_hd__nor2_1
XFILLER_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10910_ _10925_/A _10910_/B _10910_/C vssd1 vssd1 vccd1 vccd1 _10911_/A sky130_fd_sc_hd__and3_1
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11890_ _16036_/Q _11897_/C _11719_/X vssd1 vssd1 vccd1 vccd1 _11890_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ _15889_/Q _10852_/C _15034_/A vssd1 vssd1 vccd1 vccd1 _10841_/Y sky130_fd_sc_hd__a21oi_1
X_13560_ _13561_/B _13561_/C _13561_/A vssd1 vssd1 vccd1 vccd1 _13562_/B sky130_fd_sc_hd__a21o_1
X_10772_ _15878_/Q _10833_/B _10782_/C vssd1 vssd1 vccd1 vccd1 _10777_/A sky130_fd_sc_hd__and3_1
XFILLER_40_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12511_ _16123_/Q _12629_/B _12516_/C vssd1 vssd1 vccd1 vccd1 _12511_/Y sky130_fd_sc_hd__nand3_1
X_13491_ _16604_/Q vssd1 vssd1 vccd1 vccd1 _13507_/C sky130_fd_sc_hd__inv_2
XFILLER_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15230_ _15261_/C vssd1 vssd1 vccd1 vccd1 _15267_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ _16114_/Q _12493_/B _12443_/C vssd1 vssd1 vccd1 vccd1 _12442_/X sky130_fd_sc_hd__and3_1
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15161_ _16513_/Q _15267_/B _15161_/C vssd1 vssd1 vccd1 vccd1 _15169_/B sky130_fd_sc_hd__and3_1
X_12373_ _12373_/A vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__buf_2
X_14112_ _14112_/A vssd1 vssd1 vccd1 vccd1 _16349_/D sky130_fd_sc_hd__clkbuf_1
X_11324_ _11321_/Y _11330_/A _11323_/Y _11319_/C vssd1 vssd1 vccd1 vccd1 _11326_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15092_ _15090_/Y _15086_/C _15088_/Y _15089_/X vssd1 vssd1 vccd1 vccd1 _15093_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14043_ _16341_/Q _14044_/C _13986_/X vssd1 vssd1 vccd1 vccd1 _14045_/A sky130_fd_sc_hd__a21oi_1
X_11255_ _11253_/Y _11249_/C _11251_/Y _11252_/X vssd1 vssd1 vccd1 vccd1 _11256_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10206_ _15775_/Q _10402_/B _10206_/C vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__and3_1
X_11186_ _11208_/A _11186_/B _11186_/C vssd1 vssd1 vccd1 vccd1 _11187_/A sky130_fd_sc_hd__and3_1
XFILLER_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10137_ _10137_/A vssd1 vssd1 vccd1 vccd1 _15762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15994_ _16005_/CLK _15994_/D vssd1 vssd1 vccd1 vccd1 _15994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10068_ _09855_/X _10065_/B _10067_/Y vssd1 vssd1 vccd1 vccd1 _15749_/D sky130_fd_sc_hd__o21a_1
X_14945_ _15053_/A _14945_/B _14949_/B vssd1 vssd1 vccd1 vccd1 _16475_/D sky130_fd_sc_hd__nor3_1
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14876_ _14873_/Y _14874_/X _14875_/Y _14870_/C vssd1 vssd1 vccd1 vccd1 _14878_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16615_ input11/X _16615_/D vssd1 vssd1 vccd1 vccd1 _16615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13827_ _13825_/A _13825_/B _13826_/X vssd1 vssd1 vccd1 vccd1 _16308_/D sky130_fd_sc_hd__a21oi_1
XFILLER_16_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16546_ _16570_/CLK _16546_/D vssd1 vssd1 vccd1 vccd1 _16546_/Q sky130_fd_sc_hd__dfxtp_2
X_13758_ _16300_/Q _13765_/C _13698_/X vssd1 vssd1 vccd1 vccd1 _13758_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12709_ _16151_/Q _12818_/B _12718_/C vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__and3_1
X_16477_ _16607_/CLK _16477_/D vssd1 vssd1 vccd1 vccd1 _16477_/Q sky130_fd_sc_hd__dfxtp_1
X_13689_ _16291_/Q _13700_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13689_/Y sky130_fd_sc_hd__a21oi_1
X_15428_ _15440_/A vssd1 vssd1 vccd1 vccd1 _15428_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15359_ _09125_/X _15357_/A _08667_/A vssd1 vssd1 vccd1 vccd1 _15360_/B sky130_fd_sc_hd__o21ai_1
XFILLER_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09920_ _09920_/A _09920_/B vssd1 vssd1 vccd1 vccd1 _09920_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09851_ _10469_/A vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__buf_2
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _15494_/Q _08822_/C _08576_/X vssd1 vssd1 vccd1 vccd1 _08804_/B sky130_fd_sc_hd__a21oi_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09782_ _15695_/Q _09781_/C _09604_/X vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__a21o_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08733_ _08733_/A _08733_/B vssd1 vssd1 vccd1 vccd1 _08735_/A sky130_fd_sc_hd__or2_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08663_/X _08656_/A _15344_/A vssd1 vssd1 vccd1 vccd1 _08664_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ input8/X vssd1 vssd1 vccd1 vccd1 _13085_/A sky130_fd_sc_hd__buf_4
XFILLER_53_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09216_ _14911_/A vssd1 vssd1 vccd1 vccd1 _10900_/B sky130_fd_sc_hd__buf_2
XFILLER_10_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09147_ _09141_/C _09142_/C _09144_/Y _09152_/A vssd1 vssd1 vccd1 vccd1 _09152_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09078_ _09119_/A _09084_/C vssd1 vssd1 vccd1 vccd1 _09078_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08029_ _08217_/B _08029_/B vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__nand2_1
X_11040_ _15915_/Q _11212_/B _11045_/C vssd1 vssd1 vccd1 vccd1 _11040_/Y sky130_fd_sc_hd__nand3_1
XFILLER_122_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12991_ _16191_/Q _13028_/C _12933_/X vssd1 vssd1 vccd1 vccd1 _12993_/B sky130_fd_sc_hd__a21oi_1
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11942_ _16044_/Q _11950_/C _11719_/X vssd1 vssd1 vccd1 vccd1 _11942_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14730_ _14750_/C vssd1 vssd1 vccd1 vccd1 _14764_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14661_ _16432_/Q _14662_/C _14544_/X vssd1 vssd1 vccd1 vccd1 _14663_/A sky130_fd_sc_hd__a21oi_1
X_11873_ _11873_/A vssd1 vssd1 vccd1 vccd1 _16032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13612_ _13613_/B _13613_/C _13613_/A vssd1 vssd1 vccd1 vccd1 _13614_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16400_ input11/X _16400_/D vssd1 vssd1 vccd1 vccd1 _16400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10824_ _10864_/A _10824_/B _10824_/C vssd1 vssd1 vccd1 vccd1 _10825_/A sky130_fd_sc_hd__and3_1
X_14592_ _14589_/Y _14590_/X _14591_/Y _14586_/C vssd1 vssd1 vccd1 vccd1 _14594_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13543_ _13541_/A _13541_/B _13542_/X vssd1 vssd1 vccd1 vccd1 _16268_/D sky130_fd_sc_hd__a21oi_1
X_16331_ _16346_/CLK _16331_/D vssd1 vssd1 vccd1 vccd1 _16331_/Q sky130_fd_sc_hd__dfxtp_1
X_10755_ _15875_/Q _10755_/B _10755_/C vssd1 vssd1 vccd1 vccd1 _10756_/B sky130_fd_sc_hd__and3_1
X_16262_ _16533_/Q _16262_/D vssd1 vssd1 vccd1 vccd1 _16262_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13474_ _16259_/Q _13474_/B _13479_/C vssd1 vssd1 vccd1 vccd1 _13474_/Y sky130_fd_sc_hd__nand3_1
X_10686_ _10684_/Y _10685_/X _10681_/C _10682_/C vssd1 vssd1 vccd1 vccd1 _10688_/B
+ sky130_fd_sc_hd__o211ai_1
X_15213_ _15333_/A _15213_/B _15217_/B vssd1 vssd1 vccd1 vccd1 _16520_/D sky130_fd_sc_hd__nor3_1
XFILLER_139_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12425_ _16111_/Q _12462_/C _12368_/X vssd1 vssd1 vccd1 vccd1 _12427_/B sky130_fd_sc_hd__a21oi_1
X_16193_ _16555_/Q _16193_/D vssd1 vssd1 vccd1 vccd1 _16193_/Q sky130_fd_sc_hd__dfxtp_1
X_15144_ _15142_/Y _15138_/C _15140_/Y _15141_/X vssd1 vssd1 vccd1 vccd1 _15145_/C
+ sky130_fd_sc_hd__a211o_1
X_12356_ _12466_/A _12361_/C vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__or2_1
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11307_ _15954_/Q _11309_/C _11306_/X vssd1 vssd1 vccd1 vccd1 _11307_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15075_ _15180_/A _15075_/B _15079_/A vssd1 vssd1 vccd1 vccd1 _16497_/D sky130_fd_sc_hd__nor3_1
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12287_ _16092_/Q _12456_/B _12287_/C vssd1 vssd1 vccd1 vccd1 _12298_/A sky130_fd_sc_hd__and3_1
X_14026_ _14024_/Y _14020_/C _14022_/Y _14023_/X vssd1 vssd1 vccd1 vccd1 _14027_/C
+ sky130_fd_sc_hd__a211o_1
X_11238_ _12655_/A vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11169_ _11169_/A _11169_/B _11169_/C vssd1 vssd1 vccd1 vccd1 _11170_/C sky130_fd_sc_hd__or3_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15977_ _16005_/CLK _15977_/D vssd1 vssd1 vccd1 vccd1 _15977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14928_ _14936_/A _14928_/B _14928_/C vssd1 vssd1 vccd1 vccd1 _14929_/A sky130_fd_sc_hd__and3_1
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14859_ _16464_/Q _14867_/C _14858_/X vssd1 vssd1 vccd1 vccd1 _14859_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08380_ _08380_/A _08380_/B vssd1 vssd1 vccd1 vccd1 _08380_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16529_ _16595_/CLK _16529_/D vssd1 vssd1 vccd1 vccd1 _16529_/Q sky130_fd_sc_hd__dfxtp_1
X_09001_ _08832_/X _09003_/C _08924_/X vssd1 vssd1 vccd1 vccd1 _09002_/B sky130_fd_sc_hd__o21ai_1
XFILLER_144_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09903_ _09914_/C vssd1 vssd1 vccd1 vccd1 _09925_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09834_ _11269_/A vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__buf_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09765_ _09766_/B _09766_/C _09766_/A vssd1 vssd1 vccd1 vccd1 _09767_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08716_ _08721_/C vssd1 vssd1 vccd1 vccd1 _08732_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_09696_ _09691_/Y _09694_/X _09695_/Y vssd1 vssd1 vccd1 vccd1 _15674_/D sky130_fd_sc_hd__o21a_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08647_ input6/X vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__buf_4
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _15458_/Q _12932_/A _08590_/C vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__and3_1
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10540_ _10541_/B _10541_/C _10541_/A vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ _10573_/A _10471_/B vssd1 vssd1 vccd1 vccd1 _10471_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12210_ _16082_/Q _12210_/B _12212_/C vssd1 vssd1 vccd1 vccd1 _12210_/X sky130_fd_sc_hd__and3_1
XFILLER_108_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13190_ _13190_/A _13190_/B _13190_/C vssd1 vssd1 vccd1 vccd1 _13191_/A sky130_fd_sc_hd__and3_1
X_12141_ _12173_/C vssd1 vssd1 vccd1 vccd1 _12179_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_123_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12072_ _12074_/B _12074_/C _11850_/X vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__o21ai_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11023_ _13521_/A vssd1 vssd1 vccd1 vccd1 _11023_/X sky130_fd_sc_hd__clkbuf_4
X_15900_ _16553_/Q _15900_/D vssd1 vssd1 vccd1 vccd1 _15900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15831_ _16595_/CLK _15831_/D vssd1 vssd1 vccd1 vccd1 _15831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15762_ _15791_/CLK _15762_/D vssd1 vssd1 vccd1 vccd1 _15762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12974_ _16189_/Q _12975_/C _12857_/X vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__a21oi_1
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14713_ _14711_/Y _14707_/C _14709_/Y _14718_/A vssd1 vssd1 vccd1 vccd1 _14718_/B
+ sky130_fd_sc_hd__a211oi_1
X_11925_ _11940_/A _11925_/B _11925_/C vssd1 vssd1 vccd1 vccd1 _11926_/A sky130_fd_sc_hd__and3_1
X_15693_ _15791_/CLK _15693_/D vssd1 vssd1 vccd1 vccd1 _15693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11856_ _11869_/C vssd1 vssd1 vccd1 vccd1 _11878_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14644_ _14644_/A vssd1 vssd1 vccd1 vccd1 _16428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10807_ _10803_/Y _10814_/A _10806_/Y _10801_/C vssd1 vssd1 vccd1 vccd1 _10809_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14575_ _16419_/Q _14583_/C _14574_/X vssd1 vssd1 vccd1 vccd1 _14575_/Y sky130_fd_sc_hd__a21oi_1
X_11787_ _11787_/A _11787_/B vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16314_ _16346_/CLK _16314_/D vssd1 vssd1 vccd1 vccd1 _16314_/Q sky130_fd_sc_hd__dfxtp_1
X_10738_ _10738_/A _10738_/B _10738_/C vssd1 vssd1 vccd1 vccd1 _10739_/A sky130_fd_sc_hd__and3_1
X_13526_ _13526_/A _13526_/B _13526_/C vssd1 vssd1 vccd1 vccd1 _13527_/A sky130_fd_sc_hd__and3_1
XFILLER_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16245_ _16261_/CLK _16245_/D vssd1 vssd1 vccd1 vccd1 _16245_/Q sky130_fd_sc_hd__dfxtp_1
X_13457_ _16258_/Q _13459_/C _13289_/X vssd1 vssd1 vccd1 vccd1 _13457_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10669_ _15848_/Q _15847_/Q _15846_/Q _10476_/X vssd1 vssd1 vccd1 vccd1 _15858_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_127_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12408_ _16109_/Q _12409_/C _12292_/X vssd1 vssd1 vccd1 vccd1 _12410_/A sky130_fd_sc_hd__a21oi_1
X_13388_ _13388_/A _13388_/B _13388_/C vssd1 vssd1 vccd1 vccd1 _13389_/C sky130_fd_sc_hd__nand3_1
X_16176_ _16237_/CLK _16176_/D vssd1 vssd1 vccd1 vccd1 _16176_/Q sky130_fd_sc_hd__dfxtp_1
X_15127_ _15180_/A _15127_/B _15131_/A vssd1 vssd1 vccd1 vccd1 _16506_/D sky130_fd_sc_hd__nor3_1
X_12339_ _16099_/Q _12501_/B _12346_/C vssd1 vssd1 vccd1 vccd1 _12339_/X sky130_fd_sc_hd__and3_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15058_ _15058_/A vssd1 vssd1 vccd1 vccd1 _15271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14009_ _16336_/Q _14017_/C _14008_/X vssd1 vssd1 vccd1 vccd1 _14012_/B sky130_fd_sc_hd__a21o_1
XFILLER_68_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07880_ _07881_/B _08129_/A _16442_/Q vssd1 vssd1 vccd1 vccd1 _07882_/A sky130_fd_sc_hd__a21o_1
XFILLER_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16664__69 vssd1 vssd1 vccd1 vccd1 _16664__69/HI _16740_/A sky130_fd_sc_hd__conb_1
XFILLER_56_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09550_ _15648_/Q _09636_/B _09550_/C vssd1 vssd1 vccd1 vccd1 _09556_/A sky130_fd_sc_hd__and3_1
X_08501_ _08502_/A _08502_/B _08502_/C vssd1 vssd1 vccd1 vccd1 _08540_/B sky130_fd_sc_hd__a21o_1
X_09481_ _09656_/A _09481_/B vssd1 vssd1 vccd1 vccd1 _09481_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ _08410_/A _08410_/B _08431_/X vssd1 vssd1 vccd1 vccd1 _08491_/B sky130_fd_sc_hd__o21ai_1
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08363_ _08363_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _08364_/B sky130_fd_sc_hd__and2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08294_ _08294_/A _08294_/B vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__xnor2_1
XFILLER_149_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09817_ _09814_/Y _09816_/X _09809_/C _09810_/C vssd1 vssd1 vccd1 vccd1 _09819_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09748_ _09744_/X _09746_/B _09747_/Y vssd1 vssd1 vccd1 vccd1 _15684_/D sky130_fd_sc_hd__o21a_1
XFILLER_36_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _15675_/Q _09914_/B _09679_/C vssd1 vssd1 vccd1 vccd1 _09687_/A sky130_fd_sc_hd__and3_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/A vssd1 vssd1 vccd1 vccd1 _16009_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12796_/A _12690_/B _12694_/B vssd1 vssd1 vccd1 vccd1 _16147_/D sky130_fd_sc_hd__nor3_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11658_/A _11641_/B _11641_/C vssd1 vssd1 vccd1 vccd1 _11642_/A sky130_fd_sc_hd__and3_1
XFILLER_14_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _14358_/Y _14354_/C _14356_/Y _14357_/X vssd1 vssd1 vccd1 vccd1 _14361_/C
+ sky130_fd_sc_hd__a211o_1
X_11572_ _11572_/A vssd1 vssd1 vccd1 vccd1 _11586_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _16237_/Q _13364_/B _13311_/C vssd1 vssd1 vccd1 vccd1 _13319_/B sky130_fd_sc_hd__and3_1
X_10523_ _10518_/B _10521_/B _10414_/X vssd1 vssd1 vccd1 vccd1 _10524_/B sky130_fd_sc_hd__o21a_1
XFILLER_128_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ _14291_/A _14291_/B _14291_/C vssd1 vssd1 vccd1 vccd1 _14292_/C sky130_fd_sc_hd__nand3_1
X_16030_ _16118_/CLK _16030_/D vssd1 vssd1 vccd1 vccd1 _16030_/Q sky130_fd_sc_hd__dfxtp_2
X_13242_ _13242_/A vssd1 vssd1 vccd1 vccd1 _13467_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_143_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10454_ _11269_/A vssd1 vssd1 vccd1 vccd1 _10454_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ _13166_/C _13167_/C _13170_/Y _13171_/X vssd1 vssd1 vccd1 vccd1 _13174_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_123_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10385_ _10399_/A _10385_/B _10385_/C vssd1 vssd1 vccd1 vccd1 _10386_/A sky130_fd_sc_hd__and3_1
XFILLER_136_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12124_ _16069_/Q _12125_/C _12007_/X vssd1 vssd1 vccd1 vccd1 _12126_/A sky130_fd_sc_hd__a21oi_1
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12055_ _12053_/Y _12048_/C _12051_/Y _12052_/X vssd1 vssd1 vccd1 vccd1 _12056_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_77_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11006_ _11026_/C vssd1 vssd1 vccd1 vccd1 _11039_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15814_ _16595_/CLK _15814_/D vssd1 vssd1 vccd1 vccd1 _15814_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15745_ _15791_/CLK _15745_/D vssd1 vssd1 vccd1 vccd1 _15745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _16187_/Q _12967_/C _12901_/X vssd1 vssd1 vccd1 vccd1 _12957_/Y sky130_fd_sc_hd__a21oi_1
X_11908_ _11908_/A vssd1 vssd1 vccd1 vccd1 _11922_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _15791_/CLK _15676_/D vssd1 vssd1 vccd1 vccd1 _15676_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _16177_/Q _12896_/C _12887_/X vssd1 vssd1 vccd1 vccd1 _12888_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14627_ _16427_/Q _14853_/B _14633_/C vssd1 vssd1 vccd1 vccd1 _14629_/C sky130_fd_sc_hd__nand3_1
X_11839_ _11835_/Y _11845_/A _11838_/Y _11832_/C vssd1 vssd1 vccd1 vccd1 _11841_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14558_ _16403_/Q _16405_/Q _16404_/Q _10719_/X vssd1 vssd1 vccd1 vccd1 _16415_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_146_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ _13503_/C _13504_/C _13506_/Y _13507_/X vssd1 vssd1 vccd1 vccd1 _13510_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_146_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14489_ _15058_/A vssd1 vssd1 vccd1 vccd1 _14720_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_146_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16228_ _16237_/CLK _16228_/D vssd1 vssd1 vccd1 vccd1 _16228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _16261_/CLK _16159_/D vssd1 vssd1 vccd1 vccd1 _16159_/Q sky130_fd_sc_hd__dfxtp_1
X_08981_ _09142_/A _08981_/B _08981_/C vssd1 vssd1 vccd1 vccd1 _08982_/A sky130_fd_sc_hd__and3_1
XFILLER_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07932_ _07932_/A _07932_/B vssd1 vssd1 vccd1 vccd1 _07933_/B sky130_fd_sc_hd__and2_1
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07863_ _15642_/Q vssd1 vssd1 vccd1 vccd1 _09448_/C sky130_fd_sc_hd__inv_2
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ _09599_/A _09598_/Y _09599_/B vssd1 vssd1 vccd1 vccd1 _09602_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_84_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07794_ _07806_/A vssd1 vssd1 vccd1 vccd1 _07799_/A sky130_fd_sc_hd__buf_12
X_09533_ _09394_/X _09527_/B _09351_/X vssd1 vssd1 vccd1 vccd1 _09535_/A sky130_fd_sc_hd__a21oi_1
XFILLER_92_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ _15631_/Q _09472_/C _09463_/X vssd1 vssd1 vccd1 vccd1 _09468_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08415_ _08415_/A vssd1 vssd1 vccd1 vccd1 _08490_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09395_ _09394_/X _09390_/B _09351_/X vssd1 vssd1 vccd1 vccd1 _09398_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08346_ _08346_/A _08346_/B vssd1 vssd1 vccd1 vccd1 _08346_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08277_ _08092_/A _08092_/B _08276_/Y vssd1 vssd1 vccd1 vccd1 _08396_/B sky130_fd_sc_hd__o21a_1
XFILLER_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10170_ _09855_/X _10166_/B _10169_/Y vssd1 vssd1 vccd1 vccd1 _15767_/D sky130_fd_sc_hd__o21a_1
XFILLER_105_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _13860_/A vssd1 vssd1 vccd1 vccd1 _16313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12811_ _14220_/A vssd1 vssd1 vccd1 vccd1 _13377_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13791_ _13791_/A vssd1 vssd1 vccd1 vccd1 _16303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15530_ _16551_/CLK _15530_/D vssd1 vssd1 vccd1 vccd1 _15530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12740_/Y _12736_/C _12738_/Y _12747_/A vssd1 vssd1 vccd1 vccd1 _12747_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12681_/A _12673_/B _12673_/C vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__and3_1
X_15461_ _16551_/CLK _15461_/D vssd1 vssd1 vccd1 vccd1 _15461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11624_ _16571_/Q vssd1 vssd1 vccd1 vccd1 _11638_/C sky130_fd_sc_hd__inv_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _16394_/Q _14414_/C _14411_/X vssd1 vssd1 vccd1 vccd1 _14412_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15392_ _16035_/Q _16037_/Q _16036_/Q _15391_/X vssd1 vssd1 vccd1 vccd1 _16575_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_129_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11555_ _15987_/Q _11780_/B _11560_/C vssd1 vssd1 vccd1 vccd1 _11555_/Y sky130_fd_sc_hd__nand3_1
X_14343_ _16384_/Q _14351_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14347_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10506_ _10589_/A _10506_/B _10506_/C vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__and3_1
X_14274_ _14439_/A vssd1 vssd1 vccd1 vccd1 _14314_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11486_ _15979_/Q _11494_/C _11485_/X vssd1 vssd1 vccd1 vccd1 _11486_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13225_ _13246_/A _13225_/B _13225_/C vssd1 vssd1 vccd1 vccd1 _13226_/A sky130_fd_sc_hd__and3_1
X_16013_ _16554_/Q _16013_/D vssd1 vssd1 vccd1 vccd1 _16013_/Q sky130_fd_sc_hd__dfxtp_1
X_10437_ _10497_/A _10437_/B _10437_/C vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__and3_1
X_13156_ _13178_/C vssd1 vssd1 vccd1 vccd1 _13193_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _10618_/A vssd1 vssd1 vccd1 vccd1 _10573_/A sky130_fd_sc_hd__clkbuf_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12107_ _13288_/A vssd1 vssd1 vccd1 vccd1 _15247_/B sky130_fd_sc_hd__buf_2
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13087_/A _13087_/B vssd1 vssd1 vccd1 vccd1 _13093_/C sky130_fd_sc_hd__nor2_1
X_10299_ _15792_/Q _10307_/B _10138_/X vssd1 vssd1 vccd1 vccd1 _10299_/Y sky130_fd_sc_hd__a21oi_1
X_12038_ _16057_/Q _12204_/B _12038_/C vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__and3_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16634__39 vssd1 vssd1 vccd1 vccd1 _16634__39/HI _16700_/A sky130_fd_sc_hd__conb_1
XFILLER_92_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13989_ _16333_/Q _14207_/B _13989_/C vssd1 vssd1 vccd1 vccd1 _13997_/B sky130_fd_sc_hd__and3_1
X_15728_ _15812_/CLK _15728_/D vssd1 vssd1 vccd1 vccd1 _15728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15659_ _15791_/CLK _15659_/D vssd1 vssd1 vccd1 vccd1 _15659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08200_ _11113_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _08200_/X sky130_fd_sc_hd__or2_1
X_09180_ _09180_/A _09180_/B _09180_/C vssd1 vssd1 vccd1 vccd1 _09181_/C sky130_fd_sc_hd__nand3_1
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08131_ _14279_/A _07888_/B _07887_/B vssd1 vssd1 vccd1 vccd1 _08332_/A sky130_fd_sc_hd__o21ai_4
XFILLER_119_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08062_ _15633_/Q _15615_/Q vssd1 vssd1 vccd1 vccd1 _08064_/A sky130_fd_sc_hd__nand2_1
XFILLER_146_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08964_ _08923_/X _08960_/A _08924_/X vssd1 vssd1 vccd1 vccd1 _08965_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07915_ _11572_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07917_/A sky130_fd_sc_hd__or2_1
X_08895_ _15513_/Q _08896_/C _08805_/X vssd1 vssd1 vccd1 vccd1 _08898_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07846_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07846_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07777_ _07780_/A vssd1 vssd1 vccd1 vccd1 _07777_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09516_ _09514_/A _09514_/B _09513_/Y _09515_/Y vssd1 vssd1 vccd1 vccd1 _15637_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_140_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _15628_/Q _09472_/C _09252_/X vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__a21oi_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ _09378_/A _09378_/B vssd1 vssd1 vccd1 vccd1 _09378_/X sky130_fd_sc_hd__or2_1
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ _08329_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08338_/A sky130_fd_sc_hd__nand2_2
XFILLER_137_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ _11353_/C vssd1 vssd1 vccd1 vccd1 _11361_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11271_ _11267_/Y _11277_/A _11270_/Y _11264_/C vssd1 vssd1 vccd1 vccd1 _11273_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13010_ _13007_/Y _13008_/X _13009_/Y _13004_/C vssd1 vssd1 vccd1 vccd1 _13012_/B
+ sky130_fd_sc_hd__o211ai_1
X_10222_ _10322_/A _10222_/B vssd1 vssd1 vccd1 vccd1 _10222_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10153_ _15765_/Q _10308_/C _10158_/C vssd1 vssd1 vccd1 vccd1 _10153_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10084_ _10340_/A vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14961_ _14974_/C vssd1 vssd1 vccd1 vccd1 _14982_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16700_ _16700_/A _07799_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13912_ _13912_/A vssd1 vssd1 vccd1 vccd1 _16321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14892_ _14890_/A _14890_/B _14891_/X vssd1 vssd1 vccd1 vccd1 _16467_/D sky130_fd_sc_hd__a21oi_1
X_13843_ _13844_/B _13844_/C _13844_/A vssd1 vssd1 vccd1 vccd1 _13845_/B sky130_fd_sc_hd__a21o_1
XFILLER_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16562_ _16595_/CLK _16562_/D vssd1 vssd1 vccd1 vccd1 _16562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10986_ _11269_/A vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__buf_2
X_13774_ _13997_/A _13774_/B _13774_/C vssd1 vssd1 vccd1 vccd1 _13775_/C sky130_fd_sc_hd__or3_1
XFILLER_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15513_ _16551_/CLK _15513_/D vssd1 vssd1 vccd1 vccd1 _15513_/Q sky130_fd_sc_hd__dfxtp_1
X_12725_ _16154_/Q _12776_/B _12726_/C vssd1 vssd1 vccd1 vccd1 _12725_/X sky130_fd_sc_hd__and3_1
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16493_ _16607_/CLK _16493_/D vssd1 vssd1 vccd1 vccd1 _16493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15444_ _16379_/Q _16381_/Q _16380_/Q _15440_/X vssd1 vssd1 vccd1 vccd1 _16618_/D
+ sky130_fd_sc_hd__o31a_1
X_12656_ _13786_/A vssd1 vssd1 vccd1 vccd1 _12881_/B sky130_fd_sc_hd__buf_2
XFILLER_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11607_ _15996_/Q _11607_/B _11607_/C vssd1 vssd1 vccd1 vccd1 _11615_/A sky130_fd_sc_hd__and3_1
XFILLER_128_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15375_ _15933_/Q _15932_/Q _15931_/Q _15372_/X vssd1 vssd1 vccd1 vccd1 _16562_/D
+ sky130_fd_sc_hd__o31a_1
X_12587_ _12625_/A _12587_/B _12587_/C vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__and3_1
X_14326_ _14326_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14332_/C sky130_fd_sc_hd__nor2_1
X_11538_ _11536_/Y _11532_/C _11534_/Y _11535_/X vssd1 vssd1 vccd1 vccd1 _11539_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11469_ _11469_/A vssd1 vssd1 vccd1 vccd1 _15975_/D sky130_fd_sc_hd__clkbuf_1
X_14257_ _14257_/A vssd1 vssd1 vccd1 vccd1 _16370_/D sky130_fd_sc_hd__clkbuf_1
X_13208_ _14331_/A vssd1 vssd1 vccd1 vccd1 _13432_/A sky130_fd_sc_hd__clkbuf_2
X_14188_ _14184_/Y _14185_/X _14187_/Y _14182_/C vssd1 vssd1 vccd1 vccd1 _14190_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_125_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13139_ _13219_/A _13139_/B _13145_/B vssd1 vssd1 vccd1 vccd1 _16211_/D sky130_fd_sc_hd__nor3_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08680_ _08680_/A _08680_/B _08680_/C vssd1 vssd1 vccd1 vccd1 _08681_/C sky130_fd_sc_hd__nand3_1
XFILLER_39_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ _10469_/A vssd1 vssd1 vccd1 vccd1 _09301_/X sky130_fd_sc_hd__buf_2
XFILLER_34_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09232_ _09232_/A _09232_/B vssd1 vssd1 vccd1 vccd1 _09234_/A sky130_fd_sc_hd__or2_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09163_ _09294_/A vssd1 vssd1 vccd1 vccd1 _15358_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_119_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08114_ _15534_/Q _08114_/B vssd1 vssd1 vccd1 vccd1 _08114_/Y sky130_fd_sc_hd__nand2_1
X_09094_ _15557_/Q _09110_/C _09051_/X vssd1 vssd1 vccd1 vccd1 _09097_/B sky130_fd_sc_hd__a21oi_1
XFILLER_134_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08045_ _15723_/Q _15741_/Q vssd1 vssd1 vccd1 vccd1 _08046_/B sky130_fd_sc_hd__or2_1
XFILLER_135_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09996_ _09996_/A vssd1 vssd1 vccd1 vccd1 _15734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08947_ _15524_/Q _08948_/C _08777_/X vssd1 vssd1 vccd1 vccd1 _08949_/A sky130_fd_sc_hd__a21oi_1
XFILLER_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08878_ _08832_/X _08880_/C _08833_/X vssd1 vssd1 vccd1 vccd1 _08879_/B sky130_fd_sc_hd__o21ai_1
XFILLER_45_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07829_ _07830_/A vssd1 vssd1 vccd1 vccd1 _07829_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10840_ _10840_/A vssd1 vssd1 vccd1 vccd1 _15887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10771_ _15878_/Q _10812_/C _10673_/X vssd1 vssd1 vccd1 vccd1 _10773_/B sky130_fd_sc_hd__a21oi_1
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12510_ _16124_/Q _12739_/B _12510_/C vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__and3_1
X_13490_ _13490_/A vssd1 vssd1 vccd1 vccd1 _16261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12441_ _16114_/Q _12443_/C _12440_/X vssd1 vssd1 vccd1 vccd1 _12441_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15160_ _16513_/Q _15161_/C _10812_/B vssd1 vssd1 vccd1 vccd1 _15162_/A sky130_fd_sc_hd__a21oi_1
X_12372_ _16104_/Q _12380_/C _12316_/X vssd1 vssd1 vccd1 vccd1 _12376_/B sky130_fd_sc_hd__a21o_1
XFILLER_138_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11323_ _15955_/Q _11495_/B _11328_/C vssd1 vssd1 vccd1 vccd1 _11323_/Y sky130_fd_sc_hd__nand3_1
X_14111_ _14145_/A _14111_/B _14111_/C vssd1 vssd1 vccd1 vccd1 _14112_/A sky130_fd_sc_hd__and3_1
X_15091_ _15088_/Y _15089_/X _15090_/Y _15086_/C vssd1 vssd1 vccd1 vccd1 _15093_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11254_ _11251_/Y _11252_/X _11253_/Y _11249_/C vssd1 vssd1 vccd1 vccd1 _11256_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_107_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14042_ _14063_/A _14042_/B _14046_/B vssd1 vssd1 vccd1 vccd1 _16339_/D sky130_fd_sc_hd__nor3_1
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10205_ _15775_/Q _10214_/C _10204_/X vssd1 vssd1 vccd1 vccd1 _10205_/Y sky130_fd_sc_hd__a21oi_1
X_11185_ _11185_/A _11185_/B _11185_/C vssd1 vssd1 vccd1 vccd1 _11186_/C sky130_fd_sc_hd__nand3_1
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10136_ _10145_/A _10136_/B _10136_/C vssd1 vssd1 vccd1 vccd1 _10137_/A sky130_fd_sc_hd__and3_1
XFILLER_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15993_ _16005_/CLK _15993_/D vssd1 vssd1 vccd1 vccd1 _15993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10067_ _09207_/X _10065_/B _10012_/X vssd1 vssd1 vccd1 vccd1 _10067_/Y sky130_fd_sc_hd__a21oi_1
X_14944_ _14942_/Y _14936_/C _14939_/Y _14949_/A vssd1 vssd1 vccd1 vccd1 _14949_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_94_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14875_ _16465_/Q _14875_/B _14881_/C vssd1 vssd1 vccd1 vccd1 _14875_/Y sky130_fd_sc_hd__nand3_1
X_16614_ input11/X _16614_/D vssd1 vssd1 vccd1 vccd1 _16614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13826_ _13879_/A _13831_/C vssd1 vssd1 vccd1 vccd1 _13826_/X sky130_fd_sc_hd__or2_1
XFILLER_90_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16545_ _16570_/CLK _16545_/D vssd1 vssd1 vccd1 vccd1 _16545_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ _13757_/A vssd1 vssd1 vccd1 vccd1 _16298_/D sky130_fd_sc_hd__clkbuf_1
X_10969_ _15906_/Q _11076_/B _10970_/C vssd1 vssd1 vccd1 vccd1 _10969_/X sky130_fd_sc_hd__and3_1
X_12708_ _16151_/Q _12745_/C _12650_/X vssd1 vssd1 vccd1 vccd1 _12710_/B sky130_fd_sc_hd__a21oi_1
XFILLER_149_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16476_ _16607_/CLK _16476_/D vssd1 vssd1 vccd1 vccd1 _16476_/Q sky130_fd_sc_hd__dfxtp_1
X_13688_ _13688_/A vssd1 vssd1 vccd1 vccd1 _16289_/D sky130_fd_sc_hd__clkbuf_1
X_15427_ _16269_/Q _16268_/Q _16267_/Q _15422_/X vssd1 vssd1 vccd1 vccd1 _16604_/D
+ sky130_fd_sc_hd__o31a_1
X_12639_ _12637_/A _12637_/B _12638_/X vssd1 vssd1 vccd1 vccd1 _16140_/D sky130_fd_sc_hd__a21oi_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15358_ _15358_/A _15358_/B _15358_/C vssd1 vssd1 vccd1 vccd1 _15360_/A sky130_fd_sc_hd__and3_1
XFILLER_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14309_ _16379_/Q _14317_/C _14308_/X vssd1 vssd1 vccd1 vccd1 _14309_/Y sky130_fd_sc_hd__a21oi_1
X_15289_ _16707_/A _15306_/A vssd1 vssd1 vccd1 vccd1 _15291_/B sky130_fd_sc_hd__and2_1
XFILLER_144_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09850_ _09848_/A _09848_/B _09849_/X vssd1 vssd1 vccd1 vccd1 _15702_/D sky130_fd_sc_hd__a21oi_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _08807_/C vssd1 vssd1 vccd1 vccd1 _08822_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _15695_/Q _09966_/B _09781_/C vssd1 vssd1 vccd1 vccd1 _09781_/X sky130_fd_sc_hd__and3_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _15479_/Q _09271_/A _08732_/C vssd1 vssd1 vccd1 vccd1 _08733_/B sky130_fd_sc_hd__and3_1
XFILLER_38_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08663_ _10418_/A vssd1 vssd1 vccd1 vccd1 _08663_/X sky130_fd_sc_hd__buf_2
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08594_ _08594_/A vssd1 vssd1 vccd1 vccd1 _15455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09215_ input10/X vssd1 vssd1 vccd1 vccd1 _14911_/A sky130_fd_sc_hd__buf_6
XFILLER_22_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09146_ _09144_/Y _09152_/A _09141_/C _09142_/C vssd1 vssd1 vccd1 vccd1 _09148_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09077_ _09071_/B _09074_/B _08914_/X vssd1 vssd1 vccd1 vccd1 _09084_/C sky130_fd_sc_hd__o21a_1
XFILLER_135_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08028_ _08217_/A _08027_/C _15867_/Q vssd1 vssd1 vccd1 vccd1 _08029_/B sky130_fd_sc_hd__a21o_1
XFILLER_135_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ _10220_/A _09978_/X _09973_/B _08854_/A vssd1 vssd1 vccd1 vccd1 _09980_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12990_ _13022_/C vssd1 vssd1 vccd1 vccd1 _13028_/C sky130_fd_sc_hd__clkbuf_2
X_11941_ _11941_/A vssd1 vssd1 vccd1 vccd1 _16042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14660_ _14768_/A _14660_/B _14664_/B vssd1 vssd1 vccd1 vccd1 _16430_/D sky130_fd_sc_hd__nor3_1
XFILLER_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11872_ _11888_/A _11872_/B _11872_/C vssd1 vssd1 vccd1 vccd1 _11873_/A sky130_fd_sc_hd__and3_1
XFILLER_26_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13611_ _16280_/Q _13731_/B _13617_/C vssd1 vssd1 vccd1 vccd1 _13613_/C sky130_fd_sc_hd__nand3_1
X_10823_ _14954_/A _10823_/B _10823_/C vssd1 vssd1 vccd1 vccd1 _10824_/C sky130_fd_sc_hd__or3_1
XFILLER_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14591_ _16420_/Q _14591_/B _14597_/C vssd1 vssd1 vccd1 vccd1 _14591_/Y sky130_fd_sc_hd__nand3_1
X_16330_ _16346_/CLK _16330_/D vssd1 vssd1 vccd1 vccd1 _16330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ _13596_/A _13548_/C vssd1 vssd1 vccd1 vccd1 _13542_/X sky130_fd_sc_hd__or2_1
X_10754_ _15875_/Q _10755_/C _08748_/A vssd1 vssd1 vccd1 vccd1 _10756_/A sky130_fd_sc_hd__a21oi_1
XFILLER_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16261_ _16261_/CLK _16261_/D vssd1 vssd1 vccd1 vccd1 _16261_/Q sky130_fd_sc_hd__dfxtp_1
X_10685_ _15863_/Q _10735_/B _10685_/C vssd1 vssd1 vccd1 vccd1 _10685_/X sky130_fd_sc_hd__and3_1
XFILLER_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13473_ _16260_/Q _13586_/B _13473_/C vssd1 vssd1 vccd1 vccd1 _13481_/A sky130_fd_sc_hd__and3_1
X_15212_ _15210_/Y _15205_/C _15208_/Y _15217_/A vssd1 vssd1 vccd1 vccd1 _15217_/B
+ sky130_fd_sc_hd__a211oi_1
X_12424_ _12456_/C vssd1 vssd1 vccd1 vccd1 _12462_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16192_ _16555_/Q _16192_/D vssd1 vssd1 vccd1 vccd1 _16192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15143_ _15140_/Y _15141_/X _15142_/Y _15138_/C vssd1 vssd1 vccd1 vccd1 _15145_/B
+ sky130_fd_sc_hd__o211ai_1
X_12355_ _12355_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12361_/C sky130_fd_sc_hd__nor2_1
XFILLER_5_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ _13521_/A vssd1 vssd1 vccd1 vccd1 _11306_/X sky130_fd_sc_hd__buf_2
X_12286_ _16092_/Q _12296_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12286_/Y sky130_fd_sc_hd__a21oi_1
X_15074_ _16498_/Q _15074_/B _15083_/C vssd1 vssd1 vccd1 vccd1 _15079_/A sky130_fd_sc_hd__and3_1
XFILLER_113_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11237_ _15944_/Q _11246_/C _11181_/X vssd1 vssd1 vccd1 vccd1 _11242_/B sky130_fd_sc_hd__a21o_1
XFILLER_4_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14025_ _14022_/Y _14023_/X _14024_/Y _14020_/C vssd1 vssd1 vccd1 vccd1 _14027_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_141_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11168_ _11169_/B _11169_/C _10999_/X vssd1 vssd1 vccd1 vccd1 _11170_/B sky130_fd_sc_hd__o21ai_1
XFILLER_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10119_ _15777_/Q vssd1 vssd1 vccd1 vccd1 _10124_/C sky130_fd_sc_hd__inv_2
X_15976_ _16005_/CLK _15976_/D vssd1 vssd1 vccd1 vccd1 _15976_/Q sky130_fd_sc_hd__dfxtp_1
X_11099_ _15925_/Q _11099_/B _11099_/C vssd1 vssd1 vccd1 vccd1 _11109_/B sky130_fd_sc_hd__and3_1
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14927_ _14925_/Y _14921_/C _14923_/Y _14924_/X vssd1 vssd1 vccd1 vccd1 _14928_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_36_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14858_ _14858_/A vssd1 vssd1 vccd1 vccd1 _14858_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13809_ _13805_/Y _13806_/X _13808_/Y _13803_/C vssd1 vssd1 vccd1 vccd1 _13811_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14789_ _16453_/Q _14831_/C _14621_/X vssd1 vssd1 vccd1 vccd1 _14791_/B sky130_fd_sc_hd__a21oi_1
X_16528_ _16595_/CLK _16528_/D vssd1 vssd1 vccd1 vccd1 _16528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16459_ _16607_/CLK _16459_/D vssd1 vssd1 vccd1 vccd1 _16459_/Q sky130_fd_sc_hd__dfxtp_1
X_09000_ _09037_/A _09003_/C vssd1 vssd1 vccd1 vccd1 _09002_/A sky130_fd_sc_hd__and2_1
XFILLER_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09902_ _09905_/C vssd1 vssd1 vccd1 vccd1 _09914_/C sky130_fd_sc_hd__clkbuf_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _14872_/A vssd1 vssd1 vccd1 vccd1 _11269_/A sky130_fd_sc_hd__buf_4
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09764_ _15692_/Q _09867_/B _09770_/C vssd1 vssd1 vccd1 vccd1 _09766_/C sky130_fd_sc_hd__nand3_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08715_ _15489_/Q vssd1 vssd1 vccd1 vccd1 _08721_/C sky130_fd_sc_hd__inv_2
X_09695_ _09691_/Y _09694_/X _09651_/X vssd1 vssd1 vccd1 vccd1 _09695_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _08646_/A _08646_/B vssd1 vssd1 vccd1 vccd1 _15459_/D sky130_fd_sc_hd__nor2_1
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ _15458_/Q _08619_/C _08576_/X vssd1 vssd1 vccd1 vccd1 _08579_/B sky130_fd_sc_hd__a21oi_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ _10464_/B _10467_/B _10414_/X vssd1 vssd1 vccd1 vccd1 _10471_/B sky130_fd_sc_hd__o21a_1
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09129_ _15350_/A vssd1 vssd1 vccd1 vccd1 _09129_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12140_ _12160_/C vssd1 vssd1 vccd1 vccd1 _12173_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_136_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12071_ _12185_/A vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11022_ _11022_/A vssd1 vssd1 vccd1 vccd1 _15912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15830_ _16551_/CLK _15830_/D vssd1 vssd1 vccd1 vccd1 _15830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15761_ _15791_/CLK _15761_/D vssd1 vssd1 vccd1 vccd1 _15761_/Q sky130_fd_sc_hd__dfxtp_2
X_12973_ _13080_/A _12973_/B _12977_/B vssd1 vssd1 vccd1 vccd1 _16187_/D sky130_fd_sc_hd__nor3_1
XFILLER_85_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14712_ _14709_/Y _14718_/A _14711_/Y _14707_/C vssd1 vssd1 vccd1 vccd1 _14714_/B
+ sky130_fd_sc_hd__o211a_1
X_11924_ _11918_/C _11919_/C _11921_/Y _11922_/X vssd1 vssd1 vccd1 vccd1 _11925_/C
+ sky130_fd_sc_hd__a211o_1
X_15692_ _15791_/CLK _15692_/D vssd1 vssd1 vccd1 vccd1 _15692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14643_ _14651_/A _14643_/B _14643_/C vssd1 vssd1 vccd1 vccd1 _14644_/A sky130_fd_sc_hd__and3_1
X_11855_ _16575_/Q vssd1 vssd1 vccd1 vccd1 _11869_/C sky130_fd_sc_hd__clkinv_2
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _15882_/Q _10929_/B _10812_/C vssd1 vssd1 vccd1 vccd1 _10806_/Y sky130_fd_sc_hd__nand3_1
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14574_ _14858_/A vssd1 vssd1 vccd1 vccd1 _14574_/X sky130_fd_sc_hd__clkbuf_4
X_11786_ _11786_/A _11795_/B vssd1 vssd1 vccd1 vccd1 _11788_/A sky130_fd_sc_hd__or2_1
XFILLER_13_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16313_ _16346_/CLK _16313_/D vssd1 vssd1 vccd1 vccd1 _16313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _13523_/Y _13517_/C _13519_/Y _13520_/X vssd1 vssd1 vccd1 vccd1 _13526_/C
+ sky130_fd_sc_hd__a211o_1
X_10737_ _10731_/C _10732_/C _10734_/Y _10735_/X vssd1 vssd1 vccd1 vccd1 _10738_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_146_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16244_ _16261_/CLK _16244_/D vssd1 vssd1 vccd1 vccd1 _16244_/Q sky130_fd_sc_hd__dfxtp_1
X_13456_ _13456_/A vssd1 vssd1 vccd1 vccd1 _16256_/D sky130_fd_sc_hd__clkbuf_1
X_10668_ _10526_/X _10665_/B _10667_/Y vssd1 vssd1 vccd1 vccd1 _15857_/D sky130_fd_sc_hd__o21a_1
X_12407_ _12514_/A _12407_/B _12411_/B vssd1 vssd1 vccd1 vccd1 _16107_/D sky130_fd_sc_hd__nor3_1
X_16175_ _16237_/CLK _16175_/D vssd1 vssd1 vccd1 vccd1 _16175_/Q sky130_fd_sc_hd__dfxtp_1
X_13387_ _13388_/B _13388_/C _13388_/A vssd1 vssd1 vccd1 vccd1 _13389_/B sky130_fd_sc_hd__a21o_1
X_10599_ _15846_/Q _10691_/B _10606_/C vssd1 vssd1 vccd1 vccd1 _10599_/X sky130_fd_sc_hd__and3_1
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15126_ _16507_/Q _15232_/B _15135_/C vssd1 vssd1 vccd1 vccd1 _15131_/A sky130_fd_sc_hd__and3_1
X_12338_ _16099_/Q _12346_/C _12337_/X vssd1 vssd1 vccd1 vccd1 _12338_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15057_ _15057_/A _15057_/B vssd1 vssd1 vccd1 vccd1 _15059_/B sky130_fd_sc_hd__nor2_1
X_12269_ _12269_/A vssd1 vssd1 vccd1 vccd1 _12493_/B sky130_fd_sc_hd__clkbuf_2
X_14008_ _14851_/A vssd1 vssd1 vccd1 vccd1 _14008_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15959_ _15365_/A _15959_/D vssd1 vssd1 vccd1 vccd1 _15959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08500_ _08462_/A _08462_/B _08499_/Y vssd1 vssd1 vccd1 vccd1 _08502_/C sky130_fd_sc_hd__a21oi_1
X_09480_ _09655_/A _09480_/B vssd1 vssd1 vccd1 vccd1 _09481_/B sky130_fd_sc_hd__and2_1
XFILLER_64_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08431_ _08431_/A _08411_/A vssd1 vssd1 vccd1 vccd1 _08431_/X sky130_fd_sc_hd__or2b_1
XFILLER_17_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ _08363_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _08364_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08293_ _08100_/A _08100_/B _08292_/Y vssd1 vssd1 vccd1 vccd1 _08294_/B sky130_fd_sc_hd__o21a_1
XFILLER_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09816_ _15701_/Q _10190_/B _09816_/C vssd1 vssd1 vccd1 vccd1 _09816_/X sky130_fd_sc_hd__and3_1
X_09747_ _09932_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09747_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _09815_/A vssd1 vssd1 vccd1 vccd1 _09914_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08629_/A vssd1 vssd1 vccd1 vccd1 _09076_/A sky130_fd_sc_hd__buf_2
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11634_/C _11635_/C _11637_/Y _11638_/X vssd1 vssd1 vccd1 vccd1 _11641_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _11571_/A vssd1 vssd1 vccd1 vccd1 _15989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _16237_/Q _13311_/C _13140_/X vssd1 vssd1 vccd1 vccd1 _13312_/A sky130_fd_sc_hd__a21oi_1
X_10522_ _10520_/A _10520_/B _10521_/X vssd1 vssd1 vccd1 vccd1 _15828_/D sky130_fd_sc_hd__a21oi_1
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14290_ _14291_/B _14291_/C _14291_/A vssd1 vssd1 vccd1 vccd1 _14292_/B sky130_fd_sc_hd__a21o_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10453_ _10578_/A vssd1 vssd1 vccd1 vccd1 _10563_/A sky130_fd_sc_hd__clkbuf_2
X_13241_ _16227_/Q _13350_/B _13250_/C vssd1 vssd1 vccd1 vccd1 _13241_/X sky130_fd_sc_hd__and3_1
XFILLER_136_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13172_ _13170_/Y _13171_/X _13166_/C _13167_/C vssd1 vssd1 vccd1 vccd1 _13174_/B
+ sky130_fd_sc_hd__o211ai_1
X_10384_ _10384_/A _10384_/B _10384_/C vssd1 vssd1 vccd1 vccd1 _10385_/C sky130_fd_sc_hd__nand3_1
XFILLER_124_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12123_ _12230_/A _12123_/B _12127_/B vssd1 vssd1 vccd1 vccd1 _16067_/D sky130_fd_sc_hd__nor3_1
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12054_ _12051_/Y _12052_/X _12053_/Y _12048_/C vssd1 vssd1 vccd1 vccd1 _12056_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_104_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11005_ _11018_/C vssd1 vssd1 vccd1 vccd1 _11026_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15813_ _16595_/CLK _15813_/D vssd1 vssd1 vccd1 vccd1 _15813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15744_ _15791_/CLK _15744_/D vssd1 vssd1 vccd1 vccd1 _15744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12956_ _12956_/A vssd1 vssd1 vccd1 vccd1 _16185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11907_ _11907_/A vssd1 vssd1 vccd1 vccd1 _16037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _15791_/CLK _15675_/D vssd1 vssd1 vccd1 vccd1 _15675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12887_ _14015_/A vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__buf_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14911_/A vssd1 vssd1 vccd1 vccd1 _14853_/B sky130_fd_sc_hd__buf_2
X_11838_ _16027_/Q _12060_/B _11843_/C vssd1 vssd1 vccd1 vccd1 _11838_/Y sky130_fd_sc_hd__nand3_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/A vssd1 vssd1 vccd1 vccd1 _16414_/D sky130_fd_sc_hd__clkbuf_1
X_11769_ _13183_/A vssd1 vssd1 vccd1 vccd1 _12901_/A sky130_fd_sc_hd__clkbuf_4
X_13508_ _13506_/Y _13507_/X _13503_/C _13504_/C vssd1 vssd1 vccd1 vccd1 _13510_/B
+ sky130_fd_sc_hd__o211ai_1
X_14488_ _14488_/A _14488_/B vssd1 vssd1 vccd1 vccd1 _14490_/B sky130_fd_sc_hd__nor2_1
X_16227_ _16237_/CLK _16227_/D vssd1 vssd1 vccd1 vccd1 _16227_/Q sky130_fd_sc_hd__dfxtp_1
X_13439_ _16255_/Q _13479_/C _13216_/X vssd1 vssd1 vccd1 vccd1 _13442_/B sky130_fd_sc_hd__a21oi_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16158_ _16261_/CLK _16158_/D vssd1 vssd1 vccd1 vccd1 _16158_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ _16504_/Q _15267_/B _15109_/C vssd1 vssd1 vccd1 vccd1 _15117_/B sky130_fd_sc_hd__and3_1
X_08980_ _08980_/A _08980_/B _08980_/C vssd1 vssd1 vccd1 vccd1 _08981_/C sky130_fd_sc_hd__nand3_1
X_16089_ _16118_/CLK _16089_/D vssd1 vssd1 vccd1 vccd1 _16089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07931_ _07932_/A _07932_/B vssd1 vssd1 vccd1 vccd1 _07933_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07862_ _16566_/Q vssd1 vssd1 vccd1 vccd1 _11339_/A sky130_fd_sc_hd__inv_2
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09601_ _09599_/A _09599_/B _09598_/Y _09600_/Y vssd1 vssd1 vccd1 vccd1 _15655_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07793_ _07793_/A vssd1 vssd1 vccd1 vccd1 _07793_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09532_ _09529_/X _09527_/B _09531_/Y vssd1 vssd1 vccd1 vccd1 _15640_/D sky130_fd_sc_hd__o21a_1
XFILLER_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _09683_/A vssd1 vssd1 vccd1 vccd1 _09463_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08414_ _08414_/A _08414_/B vssd1 vssd1 vccd1 vccd1 _15291_/A sky130_fd_sc_hd__xor2_2
X_09394_ _09615_/A vssd1 vssd1 vccd1 vccd1 _09394_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08345_ _08345_/A _08433_/A vssd1 vssd1 vccd1 vccd1 _08407_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08276_ _16564_/Q _08276_/B vssd1 vssd1 vccd1 vccd1 _08276_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ _12810_/A vssd1 vssd1 vccd1 vccd1 _16165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13790_ _13811_/A _13790_/B _13790_/C vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__and3_1
XFILLER_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12741_ _12738_/Y _12747_/A _12740_/Y _12736_/C vssd1 vssd1 vccd1 vccd1 _12743_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _16551_/CLK _15460_/D vssd1 vssd1 vccd1 vccd1 _15460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12670_/Y _12666_/C _12668_/Y _12669_/X vssd1 vssd1 vccd1 vccd1 _12673_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14411_/A vssd1 vssd1 vccd1 vccd1 _14411_/X sky130_fd_sc_hd__buf_2
X_11623_ _11623_/A vssd1 vssd1 vccd1 vccd1 _15997_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15391_ _15409_/A vssd1 vssd1 vccd1 vccd1 _15391_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14342_ _14342_/A _14342_/B _14347_/A vssd1 vssd1 vccd1 vccd1 _16382_/D sky130_fd_sc_hd__nor3_1
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ _12686_/A vssd1 vssd1 vccd1 vccd1 _11780_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10505_ _10503_/Y _10497_/C _10500_/Y _10502_/X vssd1 vssd1 vccd1 vccd1 _10506_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14273_ _14271_/A _14271_/B _14272_/X vssd1 vssd1 vccd1 vccd1 _16372_/D sky130_fd_sc_hd__a21oi_1
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ _12968_/A vssd1 vssd1 vccd1 vccd1 _11485_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16012_ _16554_/Q _16012_/D vssd1 vssd1 vccd1 vccd1 _16012_/Q sky130_fd_sc_hd__dfxtp_1
X_13224_ _13224_/A _13224_/B _13224_/C vssd1 vssd1 vccd1 vccd1 _13225_/C sky130_fd_sc_hd__nand3_1
XFILLER_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10436_ _10436_/A _10436_/B _10436_/C vssd1 vssd1 vccd1 vccd1 _10437_/C sky130_fd_sc_hd__nand3_1
XFILLER_109_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ _13171_/C vssd1 vssd1 vccd1 vccd1 _13178_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10367_ _10365_/A _10365_/B _10366_/X vssd1 vssd1 vccd1 vccd1 _15801_/D sky130_fd_sc_hd__a21oi_1
XFILLER_112_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _16067_/Q _12218_/B _12118_/C vssd1 vssd1 vccd1 vccd1 _12106_/X sky130_fd_sc_hd__and3_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10298_/A vssd1 vssd1 vccd1 vccd1 _15789_/D sky130_fd_sc_hd__clkbuf_1
X_13086_ _14210_/A vssd1 vssd1 vccd1 vccd1 _13315_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12037_ _16057_/Q _12045_/C _12036_/X vssd1 vssd1 vccd1 vccd1 _12037_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13988_ _14830_/A vssd1 vssd1 vccd1 vccd1 _14207_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15727_ _15812_/CLK _15727_/D vssd1 vssd1 vccd1 vccd1 _15727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12939_ _16184_/Q _13164_/B _12945_/C vssd1 vssd1 vccd1 vccd1 _12941_/C sky130_fd_sc_hd__nand3_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15658_ _15791_/CLK _15658_/D vssd1 vssd1 vccd1 vccd1 _15658_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14609_ _14722_/A vssd1 vssd1 vccd1 vccd1 _14651_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15589_ _16551_/CLK _15589_/D vssd1 vssd1 vccd1 vccd1 _15589_/Q sky130_fd_sc_hd__dfxtp_2
X_08130_ _08343_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08135_/A sky130_fd_sc_hd__nor2_4
XFILLER_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08061_ _15651_/Q vssd1 vssd1 vccd1 vccd1 _09496_/C sky130_fd_sc_hd__clkinv_4
XFILLER_146_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08963_ _09124_/A _09124_/B _08963_/C vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__and3_1
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07914_ _11683_/A _07914_/B vssd1 vssd1 vccd1 vccd1 _07916_/B sky130_fd_sc_hd__xnor2_1
XFILLER_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08894_ _08946_/A _08894_/B _08898_/A vssd1 vssd1 vccd1 vccd1 _15508_/D sky130_fd_sc_hd__nor3_1
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07845_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07845_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07776_ _07780_/A vssd1 vssd1 vccd1 vccd1 _07776_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09515_ _09514_/X _09513_/Y _09424_/X vssd1 vssd1 vccd1 vccd1 _09515_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09458_/C vssd1 vssd1 vccd1 vccd1 _09472_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09377_ _09377_/A _09377_/B vssd1 vssd1 vccd1 vccd1 _09377_/Y sky130_fd_sc_hd__nor2_1
X_08328_ _08328_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08329_/A sky130_fd_sc_hd__or2_1
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08259_ _08259_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ _15947_/Q _11495_/B _11275_/C vssd1 vssd1 vccd1 vccd1 _11270_/Y sky130_fd_sc_hd__nand3_1
XFILLER_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10221_ _10215_/B _10218_/B _10164_/X vssd1 vssd1 vccd1 vccd1 _10222_/B sky130_fd_sc_hd__o21a_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10152_ _15766_/Q _10402_/B _10152_/C vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__and3_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10083_ _10083_/A vssd1 vssd1 vccd1 vccd1 _15752_/D sky130_fd_sc_hd__clkbuf_1
X_14960_ _14960_/A vssd1 vssd1 vccd1 vccd1 _14974_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13911_ _13918_/A _13911_/B _13911_/C vssd1 vssd1 vccd1 vccd1 _13912_/A sky130_fd_sc_hd__and3_1
XFILLER_101_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14891_ _15005_/A _14896_/C vssd1 vssd1 vccd1 vccd1 _14891_/X sky130_fd_sc_hd__or2_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13842_ _16312_/Q _14010_/B _13848_/C vssd1 vssd1 vccd1 vccd1 _13844_/C sky130_fd_sc_hd__nand3_1
XFILLER_47_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16561_ _16595_/CLK _16561_/D vssd1 vssd1 vccd1 vccd1 _16561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13773_ _14331_/A vssd1 vssd1 vccd1 vccd1 _13997_/A sky130_fd_sc_hd__clkbuf_2
X_10985_ _15908_/Q _11039_/B _10985_/C vssd1 vssd1 vccd1 vccd1 _10994_/A sky130_fd_sc_hd__and3_1
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15512_ _16551_/CLK _15512_/D vssd1 vssd1 vccd1 vccd1 _15512_/Q sky130_fd_sc_hd__dfxtp_1
X_12724_ _16154_/Q _12726_/C _12723_/X vssd1 vssd1 vccd1 vccd1 _12724_/Y sky130_fd_sc_hd__a21oi_1
X_16492_ _16607_/CLK _16492_/D vssd1 vssd1 vccd1 vccd1 _16492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15443_ _16373_/Q _16372_/Q _16371_/Q _15440_/X vssd1 vssd1 vccd1 vccd1 _16617_/D
+ sky130_fd_sc_hd__o31a_1
X_12655_ _12655_/A vssd1 vssd1 vccd1 vccd1 _13786_/A sky130_fd_sc_hd__buf_2
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11606_ _15996_/Q _11613_/C _11434_/X vssd1 vssd1 vccd1 vccd1 _11606_/Y sky130_fd_sc_hd__a21oi_1
X_15374_ _15925_/Q _15924_/Q _15923_/Q _15372_/X vssd1 vssd1 vccd1 vccd1 _16561_/D
+ sky130_fd_sc_hd__o31a_1
X_12586_ _12586_/A _12586_/B _12586_/C vssd1 vssd1 vccd1 vccd1 _12587_/C sky130_fd_sc_hd__or3_1
X_14325_ _14325_/A _14325_/B vssd1 vssd1 vccd1 vccd1 _14326_/B sky130_fd_sc_hd__nor2_1
X_11537_ _11534_/Y _11535_/X _11536_/Y _11532_/C vssd1 vssd1 vccd1 vccd1 _11539_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_117_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14256_ _14256_/A _14256_/B _14256_/C vssd1 vssd1 vccd1 vccd1 _14257_/A sky130_fd_sc_hd__and3_1
XFILLER_143_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11468_ _11491_/A _11468_/B _11468_/C vssd1 vssd1 vccd1 vccd1 _11469_/A sky130_fd_sc_hd__and3_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13207_ input7/X vssd1 vssd1 vccd1 vccd1 _14331_/A sky130_fd_sc_hd__clkbuf_4
X_10419_ _10418_/X _10416_/B _10224_/X vssd1 vssd1 vccd1 vccd1 _10419_/Y sky130_fd_sc_hd__a21oi_1
X_14187_ _16361_/Q _14414_/B _14187_/C vssd1 vssd1 vccd1 vccd1 _14187_/Y sky130_fd_sc_hd__nand3_1
XFILLER_124_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11399_ _11420_/C vssd1 vssd1 vccd1 vccd1 _11436_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _13136_/Y _13131_/C _13134_/Y _13145_/A vssd1 vssd1 vccd1 vccd1 _13145_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _16202_/Q _13187_/B _13076_/C vssd1 vssd1 vccd1 vccd1 _13069_/Y sky130_fd_sc_hd__nand3_1
XFILLER_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16759_ _16759_/A _07778_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09300_ _09898_/A vssd1 vssd1 vccd1 vccd1 _10469_/A sky130_fd_sc_hd__buf_2
XFILLER_62_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09231_ _15587_/Q _15346_/B _09231_/C vssd1 vssd1 vccd1 vccd1 _09232_/B sky130_fd_sc_hd__and3_1
X_09162_ _09162_/A _09162_/B vssd1 vssd1 vccd1 vccd1 _15567_/D sky130_fd_sc_hd__nor2_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08113_ _08113_/A vssd1 vssd1 vccd1 vccd1 _09016_/C sky130_fd_sc_hd__buf_2
XFILLER_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09093_ _09099_/C vssd1 vssd1 vccd1 vccd1 _09110_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08044_ _15723_/Q _15741_/Q vssd1 vssd1 vccd1 vccd1 _08046_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09995_ _10082_/A _09995_/B _09995_/C vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__and3_1
X_08946_ _08946_/A _08946_/B _08950_/B vssd1 vssd1 vccd1 vccd1 _15519_/D sky130_fd_sc_hd__nor3_1
XFILLER_88_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08877_ _09037_/A _08880_/C vssd1 vssd1 vccd1 vccd1 _08879_/A sky130_fd_sc_hd__and2_1
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07828_ _07830_/A vssd1 vssd1 vccd1 vccd1 _07828_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07759_ _07762_/A vssd1 vssd1 vccd1 vccd1 _07759_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10770_ _10805_/C vssd1 vssd1 vccd1 vccd1 _10812_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09429_ _15623_/Q _09428_/C _09383_/X vssd1 vssd1 vccd1 vccd1 _09430_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12440_ _13006_/A vssd1 vssd1 vccd1 vccd1 _12440_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12371_ _12371_/A _12371_/B _12376_/A vssd1 vssd1 vccd1 vccd1 _16102_/D sky130_fd_sc_hd__nor3_1
X_14110_ _14276_/A _14110_/B _14110_/C vssd1 vssd1 vccd1 vccd1 _14111_/C sky130_fd_sc_hd__or3_1
X_11322_ _15956_/Q _11322_/B _11322_/C vssd1 vssd1 vccd1 vccd1 _11330_/A sky130_fd_sc_hd__and3_1
XFILLER_138_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15090_ _16500_/Q _15248_/B _15090_/C vssd1 vssd1 vccd1 vccd1 _15090_/Y sky130_fd_sc_hd__nand3_1
XFILLER_126_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14041_ _14039_/Y _14035_/C _14037_/Y _14046_/A vssd1 vssd1 vccd1 vccd1 _14046_/B
+ sky130_fd_sc_hd__a211oi_1
X_11253_ _15945_/Q _11309_/B _11253_/C vssd1 vssd1 vccd1 vccd1 _11253_/Y sky130_fd_sc_hd__nand3_1
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10204_ _11269_/A vssd1 vssd1 vccd1 vccd1 _10204_/X sky130_fd_sc_hd__buf_2
XFILLER_140_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11184_ _11185_/B _11185_/C _11185_/A vssd1 vssd1 vccd1 vccd1 _11186_/B sky130_fd_sc_hd__a21o_1
XFILLER_122_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10135_ _10129_/C _10130_/C _10132_/Y _10133_/X vssd1 vssd1 vccd1 vccd1 _10136_/C
+ sky130_fd_sc_hd__a211o_1
X_15992_ _16005_/CLK _15992_/D vssd1 vssd1 vccd1 vccd1 _15992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10066_ _09851_/X _10058_/B _10062_/B _10065_/Y vssd1 vssd1 vccd1 vccd1 _15748_/D
+ sky130_fd_sc_hd__o31a_1
X_14943_ _14939_/Y _14949_/A _14942_/Y _14936_/C vssd1 vssd1 vccd1 vccd1 _14945_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14874_ _16466_/Q _15041_/B _14881_/C vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__and3_1
XFILLER_36_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13825_ _13825_/A _13825_/B vssd1 vssd1 vccd1 vccd1 _13831_/C sky130_fd_sc_hd__nor2_1
X_16613_ input11/X _16613_/D vssd1 vssd1 vccd1 vccd1 _16613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16544_ _16570_/CLK _16544_/D vssd1 vssd1 vccd1 vccd1 _16544_/Q sky130_fd_sc_hd__dfxtp_2
X_13756_ _13756_/A _13756_/B _13756_/C vssd1 vssd1 vccd1 vccd1 _13757_/A sky130_fd_sc_hd__and3_1
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10968_ _15906_/Q _10970_/C _14932_/A vssd1 vssd1 vccd1 vccd1 _10968_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _12739_/C vssd1 vssd1 vccd1 vccd1 _12745_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16475_ _16607_/CLK _16475_/D vssd1 vssd1 vccd1 vccd1 _16475_/Q sky130_fd_sc_hd__dfxtp_1
X_13687_ _13696_/A _13687_/B _13687_/C vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__and3_1
X_10899_ _15896_/Q _10907_/C _10898_/X vssd1 vssd1 vccd1 vccd1 _10902_/B sky130_fd_sc_hd__a21o_1
X_15426_ _16261_/Q _16260_/Q _16259_/Q _15422_/X vssd1 vssd1 vccd1 vccd1 _16603_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_129_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12638_ _12749_/A _12643_/C vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__or2_1
X_15357_ _15357_/A _15357_/B vssd1 vssd1 vccd1 vccd1 _16549_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12569_ _16132_/Q _12739_/B _12569_/C vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__and3_1
XFILLER_129_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14308_ _14308_/A vssd1 vssd1 vccd1 vccd1 _14308_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15288_ _15283_/C _15286_/Y _15287_/Y vssd1 vssd1 vccd1 vccd1 _16536_/D sky130_fd_sc_hd__o21a_1
XFILLER_116_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14239_ _14232_/C _14233_/C _14235_/Y _14237_/X vssd1 vssd1 vccd1 vccd1 _14240_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08800_ _15507_/Q vssd1 vssd1 vccd1 vccd1 _08807_/C sky130_fd_sc_hd__inv_2
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09780_ _09777_/A _09776_/Y _09777_/B vssd1 vssd1 vccd1 vccd1 _09780_/Y sky130_fd_sc_hd__o21bai_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _15479_/Q _08732_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _08733_/A sky130_fd_sc_hd__a21oi_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ _15274_/A vssd1 vssd1 vccd1 vccd1 _10418_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08593_ _15304_/A _08593_/B _08593_/C vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__and3_1
XFILLER_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09214_ _09256_/A _09214_/B _09222_/A vssd1 vssd1 vccd1 vccd1 _15580_/D sky130_fd_sc_hd__nor3_1
XFILLER_50_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ _15568_/Q _09145_/B _09150_/C vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__and3_1
XFILLER_108_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09076_ _09076_/A vssd1 vssd1 vccd1 vccd1 _09076_/X sky130_fd_sc_hd__buf_2
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08027_ _15867_/Q _08217_/A _08027_/C vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__nand3_1
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09978_ _14954_/A vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__buf_4
XFILLER_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08929_ _08883_/X _08926_/A _08928_/Y vssd1 vssd1 vccd1 vccd1 _15515_/D sky130_fd_sc_hd__o21a_1
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11940_ _11940_/A _11940_/B _11940_/C vssd1 vssd1 vccd1 vccd1 _11941_/A sky130_fd_sc_hd__and3_1
XFILLER_85_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11871_ _11865_/C _11866_/C _11868_/Y _11869_/X vssd1 vssd1 vccd1 vccd1 _11872_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13610_ _16280_/Q _13617_/C _13443_/X vssd1 vssd1 vccd1 vccd1 _13613_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10822_ _10823_/B _10823_/C _09978_/X vssd1 vssd1 vccd1 vccd1 _10824_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14590_ _16421_/Q _14756_/B _14597_/C vssd1 vssd1 vccd1 vccd1 _14590_/X sky130_fd_sc_hd__and3_1
XFILLER_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ _13541_/A _13541_/B vssd1 vssd1 vccd1 vccd1 _13548_/C sky130_fd_sc_hd__nor2_1
X_10753_ _10809_/A _10753_/B _10757_/B vssd1 vssd1 vccd1 vccd1 _15872_/D sky130_fd_sc_hd__nor3_1
XFILLER_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16260_ _16261_/CLK _16260_/D vssd1 vssd1 vccd1 vccd1 _16260_/Q sky130_fd_sc_hd__dfxtp_1
X_13472_ _16260_/Q _13479_/C _13414_/X vssd1 vssd1 vccd1 vccd1 _13472_/Y sky130_fd_sc_hd__a21oi_1
X_10684_ _15863_/Q _10685_/C _10492_/X vssd1 vssd1 vccd1 vccd1 _10684_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _15208_/Y _15217_/A _15210_/Y _15205_/C vssd1 vssd1 vccd1 vccd1 _15213_/B
+ sky130_fd_sc_hd__o211a_1
X_12423_ _12443_/C vssd1 vssd1 vccd1 vccd1 _12456_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16191_ _16555_/Q _16191_/D vssd1 vssd1 vccd1 vccd1 _16191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15142_ _16509_/Q _15248_/B _15142_/C vssd1 vssd1 vccd1 vccd1 _15142_/Y sky130_fd_sc_hd__nand3_1
X_12354_ _12354_/A _12354_/B vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11305_ _11305_/A vssd1 vssd1 vccd1 vccd1 _15952_/D sky130_fd_sc_hd__clkbuf_1
X_15073_ _16498_/Q _15109_/C _14906_/X vssd1 vssd1 vccd1 vccd1 _15075_/B sky130_fd_sc_hd__a21oi_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12285_ _12567_/A vssd1 vssd1 vccd1 vccd1 _12285_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14024_ _16337_/Q _14135_/B _14024_/C vssd1 vssd1 vccd1 vccd1 _14024_/Y sky130_fd_sc_hd__nand3_1
X_11236_ _11236_/A _11236_/B _11242_/A vssd1 vssd1 vccd1 vccd1 _15942_/D sky130_fd_sc_hd__nor3_1
XFILLER_106_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11167_ _11334_/A vssd1 vssd1 vccd1 vccd1 _11208_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10118_ _15749_/Q _15748_/Q _15747_/Q _09982_/X vssd1 vssd1 vccd1 vccd1 _15759_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15975_ _16005_/CLK _15975_/D vssd1 vssd1 vccd1 vccd1 _15975_/Q sky130_fd_sc_hd__dfxtp_1
X_11098_ _15925_/Q _11099_/C _10874_/X vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__a21oi_1
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10049_ _10049_/A vssd1 vssd1 vccd1 vccd1 _15745_/D sky130_fd_sc_hd__clkbuf_1
X_14926_ _14923_/Y _14924_/X _14925_/Y _14921_/C vssd1 vssd1 vccd1 vccd1 _14928_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14857_ _14857_/A vssd1 vssd1 vccd1 vccd1 _16462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _16306_/Q _14032_/B _13815_/C vssd1 vssd1 vccd1 vccd1 _13808_/Y sky130_fd_sc_hd__nand3_1
XFILLER_63_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14788_ _14823_/C vssd1 vssd1 vccd1 vccd1 _14831_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13739_ _13737_/Y _13738_/X _13733_/C _13734_/C vssd1 vssd1 vccd1 vccd1 _13741_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_32_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16527_ _16607_/CLK _16527_/D vssd1 vssd1 vccd1 vccd1 _16527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16458_ _16607_/CLK _16458_/D vssd1 vssd1 vccd1 vccd1 _16458_/Q sky130_fd_sc_hd__dfxtp_1
X_15409_ _15409_/A vssd1 vssd1 vccd1 vccd1 _15409_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16389_ _16389_/CLK _16389_/D vssd1 vssd1 vccd1 vccd1 _16389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09901_ _15596_/Q _15595_/Q _15594_/Q _09756_/X vssd1 vssd1 vccd1 vccd1 _15714_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_113_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09832_ _09832_/A vssd1 vssd1 vccd1 vccd1 _15700_/D sky130_fd_sc_hd__clkbuf_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _15692_/Q _09770_/C _09583_/X vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__a21o_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08714_ _15461_/Q _15460_/Q _15459_/Q _08667_/X vssd1 vssd1 vccd1 vccd1 _15471_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09694_ _09692_/X _09694_/B vssd1 vssd1 vccd1 vccd1 _09694_/X sky130_fd_sc_hd__and2b_1
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _08644_/X _08651_/C _15312_/A vssd1 vssd1 vccd1 vccd1 _08646_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _08843_/A vssd1 vssd1 vccd1 vccd1 _08576_/X sky130_fd_sc_hd__clkbuf_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09128_ _09128_/A _09128_/B vssd1 vssd1 vccd1 vccd1 _15559_/D sky130_fd_sc_hd__nor2_1
XFILLER_135_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09059_ _09059_/A _09059_/B _09059_/C vssd1 vssd1 vccd1 vccd1 _09060_/C sky130_fd_sc_hd__nand3_1
XFILLER_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12070_ _12068_/A _12068_/B _12069_/X vssd1 vssd1 vccd1 vccd1 _16060_/D sky130_fd_sc_hd__a21oi_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11021_ _11036_/A _11021_/B _11021_/C vssd1 vssd1 vccd1 vccd1 _11022_/A sky130_fd_sc_hd__and3_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15760_ _15791_/CLK _15760_/D vssd1 vssd1 vccd1 vccd1 _15760_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12972_ _12970_/Y _12963_/C _12966_/Y _12977_/A vssd1 vssd1 vccd1 vccd1 _12977_/B
+ sky130_fd_sc_hd__a211oi_1
X_11923_ _11921_/Y _11922_/X _11918_/C _11919_/C vssd1 vssd1 vccd1 vccd1 _11925_/B
+ sky130_fd_sc_hd__o211ai_1
X_14711_ _16439_/Q _14882_/B _14716_/C vssd1 vssd1 vccd1 vccd1 _14711_/Y sky130_fd_sc_hd__nand3_1
X_15691_ _15791_/CLK _15691_/D vssd1 vssd1 vccd1 vccd1 _15691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14642_ _14640_/Y _14636_/C _14638_/Y _14639_/X vssd1 vssd1 vccd1 vccd1 _14643_/C
+ sky130_fd_sc_hd__a211o_1
X_11854_ _11854_/A vssd1 vssd1 vccd1 vccd1 _16029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10805_ _15883_/Q _11039_/B _10805_/C vssd1 vssd1 vccd1 vccd1 _10814_/A sky130_fd_sc_hd__and3_1
X_14573_ _14573_/A vssd1 vssd1 vccd1 vccd1 _16417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11785_ _16021_/Q _11950_/B _11785_/C vssd1 vssd1 vccd1 vccd1 _11795_/B sky130_fd_sc_hd__and3_1
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16312_ _16346_/CLK _16312_/D vssd1 vssd1 vccd1 vccd1 _16312_/Q sky130_fd_sc_hd__dfxtp_1
X_13524_ _13519_/Y _13520_/X _13523_/Y _13517_/C vssd1 vssd1 vccd1 vccd1 _13526_/B
+ sky130_fd_sc_hd__o211ai_1
X_10736_ _10734_/Y _10735_/X _10731_/C _10732_/C vssd1 vssd1 vccd1 vccd1 _10738_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16243_ _16261_/CLK _16243_/D vssd1 vssd1 vccd1 vccd1 _16243_/Q sky130_fd_sc_hd__dfxtp_1
X_13455_ _13470_/A _13455_/B _13455_/C vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__and3_1
X_10667_ _09308_/X _10665_/B _10473_/X vssd1 vssd1 vccd1 vccd1 _10667_/Y sky130_fd_sc_hd__a21oi_1
X_12406_ _12404_/Y _12398_/C _12401_/Y _12411_/A vssd1 vssd1 vccd1 vccd1 _12411_/B
+ sky130_fd_sc_hd__a211oi_1
X_16174_ _16237_/CLK _16174_/D vssd1 vssd1 vccd1 vccd1 _16174_/Q sky130_fd_sc_hd__dfxtp_2
X_13386_ _16248_/Q _13445_/B _13393_/C vssd1 vssd1 vccd1 vccd1 _13388_/C sky130_fd_sc_hd__nand3_1
X_10598_ _15846_/Q _10606_/C _10393_/X vssd1 vssd1 vccd1 vccd1 _10598_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15125_ _16507_/Q _15161_/C _14906_/X vssd1 vssd1 vccd1 vccd1 _15127_/B sky130_fd_sc_hd__a21oi_1
X_12337_ _12901_/A vssd1 vssd1 vccd1 vccd1 _12337_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15056_ _15056_/A _15064_/B vssd1 vssd1 vccd1 vccd1 _15059_/A sky130_fd_sc_hd__or2_1
X_12268_ _16090_/Q _12271_/C _12157_/X vssd1 vssd1 vccd1 vccd1 _12268_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_142_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14007_ _14063_/A _14007_/B _14012_/A vssd1 vssd1 vccd1 vccd1 _16334_/D sky130_fd_sc_hd__nor3_1
X_11219_ _11219_/A _11219_/B vssd1 vssd1 vccd1 vccd1 _11220_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12199_ _12200_/B _12200_/C _12200_/A vssd1 vssd1 vccd1 vccd1 _12201_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15958_ _15365_/A _15958_/D vssd1 vssd1 vccd1 vccd1 _15958_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14909_ _14909_/A _14909_/B _14914_/A vssd1 vssd1 vccd1 vccd1 _16470_/D sky130_fd_sc_hd__nor3_1
X_15889_ _16553_/Q _15889_/D vssd1 vssd1 vccd1 vccd1 _15889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08430_ _08430_/A _08430_/B vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08361_ _08190_/A _08190_/B _08360_/X vssd1 vssd1 vccd1 vccd1 _08363_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ _15570_/Q _08292_/B vssd1 vssd1 vccd1 vccd1 _08292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09815_ _09815_/A vssd1 vssd1 vccd1 vccd1 _10190_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09746_ _09931_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09747_/B sky130_fd_sc_hd__and2_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _15675_/Q _09679_/C _09590_/X vssd1 vssd1 vccd1 vccd1 _09677_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08628_ _10307_/C vssd1 vssd1 vccd1 vccd1 _08629_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08542_/A _08542_/B _08558_/X vssd1 vssd1 vccd1 vccd1 _08567_/B sky130_fd_sc_hd__a21oi_4
XFILLER_11_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11570_ _11604_/A _11570_/B _11570_/C vssd1 vssd1 vccd1 vccd1 _11571_/A sky130_fd_sc_hd__and3_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10521_ _10521_/A _10521_/B vssd1 vssd1 vccd1 vccd1 _10521_/X sky130_fd_sc_hd__or2_1
XFILLER_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13240_ _16227_/Q _13250_/C _13184_/X vssd1 vssd1 vccd1 vccd1 _13240_/Y sky130_fd_sc_hd__a21oi_1
X_10452_ _10452_/A vssd1 vssd1 vccd1 vccd1 _15817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13171_ _16217_/Q _13336_/B _13171_/C vssd1 vssd1 vccd1 vccd1 _13171_/X sky130_fd_sc_hd__and3_1
X_10383_ _10384_/B _10384_/C _10384_/A vssd1 vssd1 vccd1 vccd1 _10385_/B sky130_fd_sc_hd__a21o_1
X_12122_ _12120_/Y _12113_/C _12117_/Y _12127_/A vssd1 vssd1 vccd1 vccd1 _12127_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_123_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12053_ _16058_/Q _12053_/B _12059_/C vssd1 vssd1 vccd1 vccd1 _12053_/Y sky130_fd_sc_hd__nand3_1
XFILLER_104_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11004_ _11004_/A vssd1 vssd1 vccd1 vccd1 _11018_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15812_ _15812_/CLK _15812_/D vssd1 vssd1 vccd1 vccd1 _15812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15743_ _15791_/CLK _15743_/D vssd1 vssd1 vccd1 vccd1 _15743_/Q sky130_fd_sc_hd__dfxtp_2
X_12955_ _12963_/A _12955_/B _12955_/C vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__and3_1
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11906_ _11940_/A _11906_/B _11906_/C vssd1 vssd1 vccd1 vccd1 _11907_/A sky130_fd_sc_hd__and3_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15791_/CLK _15674_/D vssd1 vssd1 vccd1 vccd1 _15674_/Q sky130_fd_sc_hd__dfxtp_1
X_12886_ _12886_/A vssd1 vssd1 vccd1 vccd1 _14015_/A sky130_fd_sc_hd__buf_4
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _12686_/A vssd1 vssd1 vccd1 vccd1 _12060_/B sky130_fd_sc_hd__clkbuf_2
X_14625_ _16427_/Q _14633_/C _14567_/X vssd1 vssd1 vccd1 vccd1 _14629_/B sky130_fd_sc_hd__a21o_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14556_ _14594_/A _14556_/B _14556_/C vssd1 vssd1 vccd1 vccd1 _14557_/A sky130_fd_sc_hd__and3_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11768_ _11768_/A vssd1 vssd1 vccd1 vccd1 _16017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13507_ _16265_/Q _13617_/B _13507_/C vssd1 vssd1 vccd1 vccd1 _13507_/X sky130_fd_sc_hd__and3_1
X_10719_ _14615_/A vssd1 vssd1 vccd1 vccd1 _10719_/X sky130_fd_sc_hd__buf_4
XFILLER_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ _14487_/A _14496_/B vssd1 vssd1 vccd1 vccd1 _14490_/A sky130_fd_sc_hd__or2_1
X_11699_ _11696_/Y _11698_/X _11693_/C _11694_/C vssd1 vssd1 vccd1 vccd1 _11701_/B
+ sky130_fd_sc_hd__o211ai_1
X_13438_ _13473_/C vssd1 vssd1 vccd1 vccd1 _13479_/C sky130_fd_sc_hd__clkbuf_2
X_16226_ _16237_/CLK _16226_/D vssd1 vssd1 vccd1 vccd1 _16226_/Q sky130_fd_sc_hd__dfxtp_1
X_16157_ _16555_/Q _16157_/D vssd1 vssd1 vccd1 vccd1 _16157_/Q sky130_fd_sc_hd__dfxtp_1
X_13369_ _13596_/A _13374_/C vssd1 vssd1 vccd1 vccd1 _13369_/X sky130_fd_sc_hd__or2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15108_ _16504_/Q _15109_/C _10812_/B vssd1 vssd1 vccd1 vccd1 _15110_/A sky130_fd_sc_hd__a21oi_1
XFILLER_115_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16088_ _16118_/CLK _16088_/D vssd1 vssd1 vccd1 vccd1 _16088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15039_ _15039_/A vssd1 vssd1 vccd1 vccd1 _16491_/D sky130_fd_sc_hd__clkbuf_1
X_07930_ _13435_/A _07930_/B vssd1 vssd1 vccd1 vccd1 _07932_/B sky130_fd_sc_hd__xnor2_1
XFILLER_114_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07861_ _15606_/Q vssd1 vssd1 vccd1 vccd1 _09987_/C sky130_fd_sc_hd__clkinv_2
X_09600_ _09599_/X _09598_/Y _09424_/X vssd1 vssd1 vccd1 vccd1 _09600_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07792_ _07793_/A vssd1 vssd1 vccd1 vccd1 _07792_/Y sky130_fd_sc_hd__inv_2
X_09531_ _09438_/X _09527_/B _09530_/X vssd1 vssd1 vccd1 vccd1 _09531_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09462_ _10393_/A vssd1 vssd1 vccd1 vccd1 _09683_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ _08413_/A _08428_/B vssd1 vssd1 vccd1 vccd1 _08414_/B sky130_fd_sc_hd__xnor2_2
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09393_ _09299_/X _09390_/B _09392_/Y vssd1 vssd1 vccd1 vccd1 _15613_/D sky130_fd_sc_hd__o21a_1
X_08344_ _08344_/A _08344_/B vssd1 vssd1 vccd1 vccd1 _08433_/A sky130_fd_sc_hd__xnor2_1
XFILLER_138_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08275_ _08275_/A _08275_/B vssd1 vssd1 vccd1 vccd1 _08396_/A sky130_fd_sc_hd__xnor2_4
XFILLER_138_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _09722_/C _09723_/C _09726_/Y _09733_/A vssd1 vssd1 vccd1 vccd1 _09733_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12740_ _16155_/Q _12911_/B _12745_/C vssd1 vssd1 vccd1 vccd1 _12740_/Y sky130_fd_sc_hd__nand3_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12668_/Y _12669_/X _12670_/Y _12666_/C vssd1 vssd1 vccd1 vccd1 _12673_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14410_/A vssd1 vssd1 vccd1 vccd1 _16392_/D sky130_fd_sc_hd__clkbuf_1
X_11622_ _11658_/A _11622_/B _11622_/C vssd1 vssd1 vccd1 vccd1 _11623_/A sky130_fd_sc_hd__and3_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _16027_/Q _16029_/Q _16028_/Q _15385_/X vssd1 vssd1 vccd1 vccd1 _16574_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14341_ _16383_/Q _14506_/B _14351_/C vssd1 vssd1 vccd1 vccd1 _14347_/A sky130_fd_sc_hd__and3_1
X_11553_ _15254_/B vssd1 vssd1 vccd1 vccd1 _12686_/A sky130_fd_sc_hd__buf_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10504_ _10500_/Y _10502_/X _10503_/Y _10497_/C vssd1 vssd1 vccd1 vccd1 _10506_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_7_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14272_ _14437_/A _14276_/C vssd1 vssd1 vccd1 vccd1 _14272_/X sky130_fd_sc_hd__or2_1
X_11484_ _11484_/A vssd1 vssd1 vccd1 vccd1 _15977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16011_ _16554_/Q _16011_/D vssd1 vssd1 vccd1 vccd1 _16011_/Q sky130_fd_sc_hd__dfxtp_1
X_13223_ _13224_/B _13224_/C _13224_/A vssd1 vssd1 vccd1 vccd1 _13225_/B sky130_fd_sc_hd__a21o_1
X_10435_ _10436_/B _10436_/C _10436_/A vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__a21o_1
XFILLER_124_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13154_ _16598_/Q vssd1 vssd1 vccd1 vccd1 _13171_/C sky130_fd_sc_hd__inv_2
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10366_ _10521_/A _10366_/B vssd1 vssd1 vccd1 vccd1 _10366_/X sky130_fd_sc_hd__or2_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _16067_/Q _12118_/C _12050_/X vssd1 vssd1 vccd1 vccd1 _12105_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13085_ _13085_/A vssd1 vssd1 vccd1 vccd1 _14210_/A sky130_fd_sc_hd__clkbuf_4
X_10297_ _10338_/A _10297_/B _10297_/C vssd1 vssd1 vccd1 vccd1 _10298_/A sky130_fd_sc_hd__and3_1
XFILLER_105_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12036_ _12605_/A vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13987_ _16333_/Q _13989_/C _13986_/X vssd1 vssd1 vccd1 vccd1 _13990_/A sky130_fd_sc_hd__a21oi_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15726_ _16551_/CLK _15726_/D vssd1 vssd1 vccd1 vccd1 _15726_/Q sky130_fd_sc_hd__dfxtp_2
X_12938_ _13786_/A vssd1 vssd1 vccd1 vccd1 _13164_/B sky130_fd_sc_hd__clkbuf_4
X_15657_ _15791_/CLK _15657_/D vssd1 vssd1 vccd1 vccd1 _15657_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12869_ _12907_/A _12869_/B _12869_/C vssd1 vssd1 vccd1 vccd1 _12870_/A sky130_fd_sc_hd__and3_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ _14606_/A _14606_/B _14607_/X vssd1 vssd1 vccd1 vccd1 _16422_/D sky130_fd_sc_hd__a21oi_1
XFILLER_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15588_ _16570_/CLK _15588_/D vssd1 vssd1 vccd1 vccd1 _15588_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14539_ _16413_/Q _14710_/B _14539_/C vssd1 vssd1 vccd1 vccd1 _14549_/A sky130_fd_sc_hd__and3_1
XFILLER_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08060_ _16469_/Q vssd1 vssd1 vccd1 vccd1 _14785_/A sky130_fd_sc_hd__clkinv_2
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16209_ _16237_/CLK _16209_/D vssd1 vssd1 vccd1 vccd1 _16209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08962_ _10414_/A vssd1 vssd1 vccd1 vccd1 _09124_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07913_ _13212_/A _08151_/B vssd1 vssd1 vccd1 vccd1 _07914_/B sky130_fd_sc_hd__xnor2_4
X_08893_ _15512_/Q _09053_/B _08896_/C vssd1 vssd1 vccd1 vccd1 _08898_/A sky130_fd_sc_hd__and3_1
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07844_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07844_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07775_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07780_/A sky130_fd_sc_hd__buf_12
X_09514_ _09514_/A _09514_/B vssd1 vssd1 vccd1 vccd1 _09514_/X sky130_fd_sc_hd__or2_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09445_ _09448_/C vssd1 vssd1 vccd1 vccd1 _09458_/C sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _15613_/Q _09837_/A _09382_/C vssd1 vssd1 vccd1 vccd1 _09378_/B sky130_fd_sc_hd__and3_1
X_08327_ _08327_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08339_/A sky130_fd_sc_hd__nand2_2
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08258_ _08259_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _08458_/A sky130_fd_sc_hd__or2_4
XFILLER_119_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08189_ _08360_/B _08189_/B vssd1 vssd1 vccd1 vccd1 _08190_/B sky130_fd_sc_hd__xnor2_2
XFILLER_106_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10220_ _10220_/A vssd1 vssd1 vccd1 vccd1 _10220_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _14941_/A vssd1 vssd1 vccd1 vccd1 _10402_/B sky130_fd_sc_hd__clkbuf_2
X_10082_ _10082_/A _10082_/B _10082_/C vssd1 vssd1 vccd1 vccd1 _10083_/A sky130_fd_sc_hd__and3_1
XFILLER_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13910_ _13908_/Y _13903_/C _13905_/Y _13906_/X vssd1 vssd1 vccd1 vccd1 _13911_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14890_ _14890_/A _14890_/B vssd1 vssd1 vccd1 vccd1 _14896_/C sky130_fd_sc_hd__nor2_1
X_13841_ _16312_/Q _13848_/C _13729_/X vssd1 vssd1 vccd1 vccd1 _13844_/B sky130_fd_sc_hd__a21o_1
XFILLER_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16560_ _16595_/CLK _16560_/D vssd1 vssd1 vccd1 vccd1 _16560_/Q sky130_fd_sc_hd__dfxtp_1
X_13772_ _13774_/B _13774_/C _13546_/X vssd1 vssd1 vccd1 vccd1 _13775_/B sky130_fd_sc_hd__o21ai_1
XFILLER_16_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10984_ _15908_/Q _10992_/C _10866_/X vssd1 vssd1 vccd1 vccd1 _10984_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15511_ _16551_/CLK _15511_/D vssd1 vssd1 vccd1 vccd1 _15511_/Q sky130_fd_sc_hd__dfxtp_2
X_12723_ _13006_/A vssd1 vssd1 vccd1 vccd1 _12723_/X sky130_fd_sc_hd__buf_2
X_16491_ _16607_/CLK _16491_/D vssd1 vssd1 vccd1 vccd1 _16491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12654_ _16144_/Q _12663_/C _12598_/X vssd1 vssd1 vccd1 vccd1 _12659_/B sky130_fd_sc_hd__a21o_1
X_15442_ _16363_/Q _16365_/Q _16364_/Q _15440_/X vssd1 vssd1 vccd1 vccd1 _16616_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_130_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _11605_/A vssd1 vssd1 vccd1 vccd1 _15994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15373_ _15917_/Q _15916_/Q _15915_/Q _15372_/X vssd1 vssd1 vccd1 vccd1 _16560_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_128_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12585_ _12586_/B _12586_/C _12416_/X vssd1 vssd1 vccd1 vccd1 _12587_/B sky130_fd_sc_hd__o21ai_1
X_11536_ _15985_/Q _11594_/B _11536_/C vssd1 vssd1 vccd1 vccd1 _11536_/Y sky130_fd_sc_hd__nand3_1
X_14324_ _14324_/A _14332_/B vssd1 vssd1 vccd1 vccd1 _14326_/A sky130_fd_sc_hd__or2_1
XFILLER_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14255_ _14253_/Y _14248_/C _14250_/Y _14252_/X vssd1 vssd1 vccd1 vccd1 _14256_/C
+ sky130_fd_sc_hd__a211o_1
X_11467_ _11467_/A _11467_/B _11467_/C vssd1 vssd1 vccd1 vccd1 _11468_/C sky130_fd_sc_hd__nand3_1
XFILLER_137_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13206_ _13209_/B _13209_/C _12982_/X vssd1 vssd1 vccd1 vccd1 _13210_/B sky130_fd_sc_hd__o21ai_1
XFILLER_143_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10418_ _10418_/A vssd1 vssd1 vccd1 vccd1 _10418_/X sky130_fd_sc_hd__clkbuf_2
X_14186_ _14186_/A vssd1 vssd1 vccd1 vccd1 _14414_/B sky130_fd_sc_hd__clkbuf_2
X_11398_ _11412_/C vssd1 vssd1 vccd1 vccd1 _11420_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13137_ _13134_/Y _13145_/A _13136_/Y _13131_/C vssd1 vssd1 vccd1 vccd1 _13139_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _15800_/Q _10396_/B _10355_/C vssd1 vssd1 vccd1 vccd1 _10349_/Y sky130_fd_sc_hd__nand3_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13068_ _16203_/Q _13068_/B _13076_/C vssd1 vssd1 vccd1 vccd1 _13068_/X sky130_fd_sc_hd__and3_1
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12019_ _12056_/A _12019_/B _12019_/C vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__and3_1
XFILLER_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16758_ _16758_/A _07777_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
XFILLER_81_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15709_ _15812_/CLK _15709_/D vssd1 vssd1 vccd1 vccd1 _15709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16689_ _16689_/A _07786_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_110_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09230_ _15587_/Q _09231_/C _10510_/A vssd1 vssd1 vccd1 vccd1 _09232_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ _09038_/X _09165_/C _09126_/X vssd1 vssd1 vccd1 vccd1 _09162_/B sky130_fd_sc_hd__o21ai_1
XFILLER_119_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08112_ _07855_/A _08106_/B _08111_/X vssd1 vssd1 vccd1 vccd1 _08306_/A sky130_fd_sc_hd__o21ai_2
XFILLER_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09092_ _15570_/Q vssd1 vssd1 vccd1 vccd1 _09099_/C sky130_fd_sc_hd__inv_2
XFILLER_119_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ _15759_/Q vssd1 vssd1 vccd1 vccd1 _10029_/C sky130_fd_sc_hd__inv_2
XFILLER_115_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09994_ _09994_/A _09994_/B _09994_/C vssd1 vssd1 vccd1 vccd1 _09995_/C sky130_fd_sc_hd__nand3_1
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08945_ _08939_/C _08940_/C _08942_/Y _08950_/A vssd1 vssd1 vccd1 vccd1 _08950_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08876_ _10016_/A vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07827_ _07830_/A vssd1 vssd1 vccd1 vccd1 _07827_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07758_ _07762_/A vssd1 vssd1 vccd1 vccd1 _07758_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09428_ _15623_/Q _09472_/B _09428_/C vssd1 vssd1 vccd1 vccd1 _09428_/X sky130_fd_sc_hd__and3_1
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09359_ _15610_/Q _09382_/C _09252_/X vssd1 vssd1 vccd1 vccd1 _09361_/B sky130_fd_sc_hd__a21oi_1
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12370_ _16103_/Q _12535_/B _12380_/C vssd1 vssd1 vccd1 vccd1 _12376_/A sky130_fd_sc_hd__and3_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11321_ _15956_/Q _11328_/C _11150_/X vssd1 vssd1 vccd1 vccd1 _11321_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14040_ _14037_/Y _14046_/A _14039_/Y _14035_/C vssd1 vssd1 vccd1 vccd1 _14042_/B
+ sky130_fd_sc_hd__o211a_1
X_11252_ _15946_/Q _11359_/B _11253_/C vssd1 vssd1 vccd1 vccd1 _11252_/X sky130_fd_sc_hd__and3_1
X_10203_ _10578_/A vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ _15936_/Q _11183_/B _11190_/C vssd1 vssd1 vccd1 vccd1 _11185_/C sky130_fd_sc_hd__nand3_1
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10134_ _10132_/Y _10133_/X _10129_/C _10130_/C vssd1 vssd1 vccd1 vccd1 _10136_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_95_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15991_ _16005_/CLK _15991_/D vssd1 vssd1 vccd1 vccd1 _15991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10065_ _10065_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _10065_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14942_ _16475_/Q _15156_/B _14947_/C vssd1 vssd1 vccd1 vccd1 _14942_/Y sky130_fd_sc_hd__nand3_1
XFILLER_125_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14873_ _16466_/Q _14881_/C _14872_/X vssd1 vssd1 vccd1 vccd1 _14873_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16612_ input11/X _16612_/D vssd1 vssd1 vccd1 vccd1 _16612_/Q sky130_fd_sc_hd__dfxtp_1
X_13824_ _13824_/A _13824_/B vssd1 vssd1 vccd1 vccd1 _13825_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16543_ _16570_/CLK _16543_/D vssd1 vssd1 vccd1 vccd1 _16703_/A sky130_fd_sc_hd__dfxtp_2
X_10967_ _10967_/A vssd1 vssd1 vccd1 vccd1 _15904_/D sky130_fd_sc_hd__clkbuf_1
X_13755_ _13753_/Y _13748_/C _13751_/Y _13752_/X vssd1 vssd1 vccd1 vccd1 _13756_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12706_ _12726_/C vssd1 vssd1 vccd1 vccd1 _12739_/C sky130_fd_sc_hd__clkbuf_1
X_16474_ _16607_/CLK _16474_/D vssd1 vssd1 vccd1 vccd1 _16474_/Q sky130_fd_sc_hd__dfxtp_1
X_10898_ _12029_/A vssd1 vssd1 vccd1 vccd1 _10898_/X sky130_fd_sc_hd__buf_2
X_13686_ _13684_/Y _13679_/C _13681_/Y _13683_/X vssd1 vssd1 vccd1 vccd1 _13687_/C
+ sky130_fd_sc_hd__a211o_1
X_15425_ _16253_/Q _16252_/Q _16251_/Q _15422_/X vssd1 vssd1 vccd1 vccd1 _16602_/D
+ sky130_fd_sc_hd__o31a_1
X_12637_ _12637_/A _12637_/B vssd1 vssd1 vccd1 vccd1 _12643_/C sky130_fd_sc_hd__nor2_1
XFILLER_129_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15356_ _09744_/A _15358_/C _08667_/A vssd1 vssd1 vccd1 vccd1 _15357_/B sky130_fd_sc_hd__o21ai_1
X_12568_ _16132_/Q _12578_/C _12567_/X vssd1 vssd1 vccd1 vccd1 _12568_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11519_ _15983_/Q _11688_/B _11529_/C vssd1 vssd1 vccd1 vccd1 _11525_/A sky130_fd_sc_hd__and3_1
X_14307_ _14307_/A vssd1 vssd1 vccd1 vccd1 _16377_/D sky130_fd_sc_hd__clkbuf_1
X_15287_ _15283_/C _15286_/Y _10716_/X vssd1 vssd1 vccd1 vccd1 _15287_/Y sky130_fd_sc_hd__a21oi_1
X_12499_ _12499_/A vssd1 vssd1 vccd1 vccd1 _16121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14238_ _14235_/Y _14237_/X _14232_/C _14233_/C vssd1 vssd1 vccd1 vccd1 _14240_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14169_ _16359_/Q _14207_/C _14060_/X vssd1 vssd1 vccd1 vccd1 _14171_/B sky130_fd_sc_hd__a21oi_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _08730_/A _08730_/B _08734_/B vssd1 vssd1 vccd1 vccd1 _15474_/D sky130_fd_sc_hd__nor3_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08661_ _10276_/A vssd1 vssd1 vccd1 vccd1 _08661_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08592_ _08592_/A _08592_/B _08592_/C vssd1 vssd1 vccd1 vccd1 _08593_/C sky130_fd_sc_hd__nand3_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ _15584_/Q _15332_/B _09220_/C vssd1 vssd1 vccd1 vccd1 _09222_/A sky130_fd_sc_hd__and3_1
XFILLER_139_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09144_ _15568_/Q _09150_/C _09063_/X vssd1 vssd1 vccd1 vccd1 _09144_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09075_ _09073_/A _09073_/B _09074_/X vssd1 vssd1 vccd1 vccd1 _15547_/D sky130_fd_sc_hd__a21oi_1
X_08026_ _15849_/Q _15831_/Q vssd1 vssd1 vccd1 vccd1 _08027_/C sky130_fd_sc_hd__or2_1
XFILLER_116_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09977_ _08654_/X _09973_/B _09792_/X vssd1 vssd1 vccd1 vccd1 _09980_/A sky130_fd_sc_hd__a21oi_1
XFILLER_104_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08928_ _08796_/X _08926_/A _08927_/X vssd1 vssd1 vccd1 vccd1 _08928_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08859_ _10447_/A vssd1 vssd1 vccd1 vccd1 _08859_/X sky130_fd_sc_hd__buf_2
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11870_ _11868_/Y _11869_/X _11865_/C _11866_/C vssd1 vssd1 vccd1 vccd1 _11872_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_26_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10821_ _11051_/A vssd1 vssd1 vccd1 vccd1 _10864_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ _10750_/Y _10746_/C _10748_/Y _10757_/A vssd1 vssd1 vccd1 vccd1 _10757_/B
+ sky130_fd_sc_hd__a211oi_1
X_13540_ _13540_/A _13540_/B vssd1 vssd1 vccd1 vccd1 _13541_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ _13471_/A vssd1 vssd1 vccd1 vccd1 _16258_/D sky130_fd_sc_hd__clkbuf_1
X_10683_ _10683_/A vssd1 vssd1 vccd1 vccd1 _15860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15210_ _16520_/Q _15262_/B _15215_/C vssd1 vssd1 vccd1 vccd1 _15210_/Y sky130_fd_sc_hd__nand3_1
X_12422_ _12435_/C vssd1 vssd1 vccd1 vccd1 _12443_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16190_ _16555_/Q _16190_/D vssd1 vssd1 vccd1 vccd1 _16190_/Q sky130_fd_sc_hd__dfxtp_2
X_15141_ _16510_/Q _15247_/B _15142_/C vssd1 vssd1 vccd1 vccd1 _15141_/X sky130_fd_sc_hd__and3_1
X_12353_ _12353_/A _12361_/B vssd1 vssd1 vccd1 vccd1 _12355_/A sky130_fd_sc_hd__or2_1
XFILLER_126_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11304_ _11319_/A _11304_/B _11304_/C vssd1 vssd1 vccd1 vccd1 _11305_/A sky130_fd_sc_hd__and3_1
X_15072_ _15103_/C vssd1 vssd1 vccd1 vccd1 _15109_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_107_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12284_ _12284_/A vssd1 vssd1 vccd1 vccd1 _16090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14023_ _16338_/Q _14185_/B _14024_/C vssd1 vssd1 vccd1 vccd1 _14023_/X sky130_fd_sc_hd__and3_1
X_11235_ _15943_/Q _11402_/B _11246_/C vssd1 vssd1 vccd1 vccd1 _11242_/A sky130_fd_sc_hd__and3_1
XFILLER_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11166_ _11164_/A _11164_/B _11165_/X vssd1 vssd1 vccd1 vccd1 _15932_/D sky130_fd_sc_hd__a21oi_1
XFILLER_68_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10117_ _09855_/X _10114_/B _10116_/Y vssd1 vssd1 vccd1 vccd1 _15758_/D sky130_fd_sc_hd__o21a_1
XFILLER_121_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15974_ _16005_/CLK _15974_/D vssd1 vssd1 vccd1 vccd1 _15974_/Q sky130_fd_sc_hd__dfxtp_2
X_11097_ _11097_/A _11097_/B _11101_/B vssd1 vssd1 vccd1 vccd1 _15923_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10048_ _10082_/A _10048_/B _10048_/C vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__and3_1
X_14925_ _16473_/Q _14982_/B _14925_/C vssd1 vssd1 vccd1 vccd1 _14925_/Y sky130_fd_sc_hd__nand3_1
XFILLER_75_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14856_ _14878_/A _14856_/B _14856_/C vssd1 vssd1 vccd1 vccd1 _14857_/A sky130_fd_sc_hd__and3_1
XFILLER_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13807_ _14647_/A vssd1 vssd1 vccd1 vccd1 _14032_/B sky130_fd_sc_hd__clkbuf_2
X_14787_ _14808_/C vssd1 vssd1 vccd1 vccd1 _14823_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11999_ _11999_/A vssd1 vssd1 vccd1 vccd1 _16050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16526_ _16595_/CLK _16526_/D vssd1 vssd1 vccd1 vccd1 _16526_/Q sky130_fd_sc_hd__dfxtp_1
X_13738_ _16297_/Q _13900_/B _13738_/C vssd1 vssd1 vccd1 vccd1 _13738_/X sky130_fd_sc_hd__and3_1
XFILLER_32_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16457_ _16607_/CLK _16457_/D vssd1 vssd1 vccd1 vccd1 _16457_/Q sky130_fd_sc_hd__dfxtp_1
X_13669_ _13670_/B _13670_/C _13670_/A vssd1 vssd1 vccd1 vccd1 _13671_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15408_ _16149_/Q _16148_/Q _16147_/Q _15403_/X vssd1 vssd1 vccd1 vccd1 _16589_/D
+ sky130_fd_sc_hd__o31a_1
X_16388_ _16389_/CLK _16388_/D vssd1 vssd1 vccd1 vccd1 _16388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15339_ _15339_/A vssd1 vssd1 vccd1 vccd1 _16545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _15713_/D sky130_fd_sc_hd__nor2_1
XFILLER_144_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09831_ _09951_/A _09831_/B _09831_/C vssd1 vssd1 vccd1 vccd1 _09832_/A sky130_fd_sc_hd__and3_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09841_/A _09762_/B _09766_/A vssd1 vssd1 vccd1 vccd1 _15688_/D sky130_fd_sc_hd__nor3_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16675__80 vssd1 vssd1 vccd1 vccd1 _16675__80/HI _16751_/A sky130_fd_sc_hd__conb_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08661_/X _08710_/A _08712_/Y vssd1 vssd1 vccd1 vccd1 _15470_/D sky130_fd_sc_hd__o21a_1
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09693_ _15677_/Q _09692_/C _09604_/X vssd1 vssd1 vccd1 vccd1 _09694_/B sky130_fd_sc_hd__a21o_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08644_ _09038_/A vssd1 vssd1 vccd1 vccd1 _08644_/X sky130_fd_sc_hd__buf_2
XFILLER_94_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08575_ _14906_/A vssd1 vssd1 vccd1 vccd1 _08843_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09127_ _09125_/X _09123_/A _09126_/X vssd1 vssd1 vccd1 vccd1 _09128_/B sky130_fd_sc_hd__o21ai_1
XFILLER_148_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ _09059_/B _09059_/C _09059_/A vssd1 vssd1 vccd1 vccd1 _09060_/B sky130_fd_sc_hd__a21o_1
XFILLER_136_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08009_ _16619_/Q vssd1 vssd1 vccd1 vccd1 _14335_/A sky130_fd_sc_hd__clkinv_4
XFILLER_150_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11020_ _11014_/C _11015_/C _11017_/Y _11018_/X vssd1 vssd1 vccd1 vccd1 _11021_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12971_ _12966_/Y _12977_/A _12970_/Y _12963_/C vssd1 vssd1 vccd1 vccd1 _12973_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14710_ _16440_/Q _14710_/B _14710_/C vssd1 vssd1 vccd1 vccd1 _14718_/A sky130_fd_sc_hd__and3_1
X_11922_ _16041_/Q _11922_/B _11922_/C vssd1 vssd1 vccd1 vccd1 _11922_/X sky130_fd_sc_hd__and3_1
X_15690_ _15791_/CLK _15690_/D vssd1 vssd1 vccd1 vccd1 _15690_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14641_ _14638_/Y _14639_/X _14640_/Y _14636_/C vssd1 vssd1 vccd1 vccd1 _14643_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11853_ _11888_/A _11853_/B _11853_/C vssd1 vssd1 vccd1 vccd1 _11854_/A sky130_fd_sc_hd__and3_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10804_ _14821_/A vssd1 vssd1 vccd1 vccd1 _11039_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11784_ _16021_/Q _11785_/C _11726_/X vssd1 vssd1 vccd1 vccd1 _11786_/A sky130_fd_sc_hd__a21oi_1
X_14572_ _14594_/A _14572_/B _14572_/C vssd1 vssd1 vccd1 vccd1 _14573_/A sky130_fd_sc_hd__and3_1
X_16311_ _16346_/CLK _16311_/D vssd1 vssd1 vccd1 vccd1 _16311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _16266_/Q _13753_/B _13531_/C vssd1 vssd1 vccd1 vccd1 _13523_/Y sky130_fd_sc_hd__nand3_1
X_10735_ _15872_/Q _10735_/B _10735_/C vssd1 vssd1 vccd1 vccd1 _10735_/X sky130_fd_sc_hd__and3_1
XFILLER_9_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16242_ _16261_/CLK _16242_/D vssd1 vssd1 vccd1 vccd1 _16242_/Q sky130_fd_sc_hd__dfxtp_1
X_13454_ _13447_/C _13448_/C _13451_/Y _13452_/X vssd1 vssd1 vccd1 vccd1 _13455_/C
+ sky130_fd_sc_hd__a211o_1
X_10666_ _10469_/X _10659_/B _10662_/B _10665_/Y vssd1 vssd1 vccd1 vccd1 _15856_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12405_ _12401_/Y _12411_/A _12404_/Y _12398_/C vssd1 vssd1 vccd1 vccd1 _12407_/B
+ sky130_fd_sc_hd__o211a_1
X_13385_ _16248_/Q _13393_/C _13162_/X vssd1 vssd1 vccd1 vccd1 _13388_/B sky130_fd_sc_hd__a21o_1
X_16173_ _16555_/Q _16173_/D vssd1 vssd1 vccd1 vccd1 _16173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10597_ _10597_/A vssd1 vssd1 vccd1 vccd1 _15843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ _15155_/C vssd1 vssd1 vccd1 vccd1 _15161_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12336_ _12336_/A vssd1 vssd1 vccd1 vccd1 _16097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15055_ _16495_/Q _15055_/B _15055_/C vssd1 vssd1 vccd1 vccd1 _15064_/B sky130_fd_sc_hd__and3_1
X_12267_ _12267_/A vssd1 vssd1 vccd1 vccd1 _16088_/D sky130_fd_sc_hd__clkbuf_1
X_11218_ _11218_/A _11226_/B vssd1 vssd1 vccd1 vccd1 _11220_/A sky130_fd_sc_hd__or2_1
X_14006_ _16335_/Q _14227_/B _14017_/C vssd1 vssd1 vccd1 vccd1 _14012_/A sky130_fd_sc_hd__and3_1
X_12198_ _16080_/Q _12318_/B _12204_/C vssd1 vssd1 vccd1 vccd1 _12200_/C sky130_fd_sc_hd__nand3_1
XFILLER_122_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11149_ _11149_/A vssd1 vssd1 vccd1 vccd1 _15930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15957_ _16005_/CLK _15957_/D vssd1 vssd1 vccd1 vccd1 _15957_/Q sky130_fd_sc_hd__dfxtp_1
X_14908_ _16471_/Q _15074_/B _14918_/C vssd1 vssd1 vccd1 vccd1 _14914_/A sky130_fd_sc_hd__and3_1
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15888_ _16553_/Q _15888_/D vssd1 vssd1 vccd1 vccd1 _15888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14839_ _14839_/A _14839_/B _14839_/C vssd1 vssd1 vccd1 vccd1 _14840_/C sky130_fd_sc_hd__or3_1
X_08360_ _08189_/B _08360_/B vssd1 vssd1 vccd1 vccd1 _08360_/X sky130_fd_sc_hd__and2b_1
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16509_ _16607_/CLK _16509_/D vssd1 vssd1 vccd1 vccd1 _16509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08291_ _08291_/A _08291_/B vssd1 vssd1 vccd1 vccd1 _08294_/A sky130_fd_sc_hd__xnor2_1
XFILLER_149_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09814_ _15701_/Q _09816_/C _09813_/X vssd1 vssd1 vccd1 vccd1 _09814_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09745_ _09737_/Y _09739_/X _09741_/B vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__o21a_1
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09676_/A vssd1 vssd1 vccd1 vccd1 _15671_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _10456_/A vssd1 vssd1 vccd1 vccd1 _10307_/C sky130_fd_sc_hd__buf_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _08543_/A _08543_/B _08541_/A vssd1 vssd1 vccd1 vccd1 _08558_/X sky130_fd_sc_hd__a21o_1
X_08489_ _08489_/A vssd1 vssd1 vccd1 vccd1 _15449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10520_ _10520_/A _10520_/B vssd1 vssd1 vccd1 vccd1 _10521_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _10497_/A _10451_/B _10451_/C vssd1 vssd1 vccd1 vccd1 _10452_/A sky130_fd_sc_hd__and3_1
X_13170_ _16217_/Q _13178_/C _13169_/X vssd1 vssd1 vccd1 vccd1 _13170_/Y sky130_fd_sc_hd__a21oi_1
X_10382_ _15808_/Q _10434_/B _10388_/C vssd1 vssd1 vccd1 vccd1 _10384_/C sky130_fd_sc_hd__nand3_1
XFILLER_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12121_ _12117_/Y _12127_/A _12120_/Y _12113_/C vssd1 vssd1 vccd1 vccd1 _12123_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12052_ _16059_/Q _12218_/B _12059_/C vssd1 vssd1 vccd1 vccd1 _12052_/X sky130_fd_sc_hd__and3_1
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11003_ _11003_/A vssd1 vssd1 vccd1 vccd1 _15909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15811_ _15812_/CLK _15811_/D vssd1 vssd1 vccd1 vccd1 _15811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15742_ _15791_/CLK _15742_/D vssd1 vssd1 vccd1 vccd1 _15742_/Q sky130_fd_sc_hd__dfxtp_2
X_12954_ _12952_/Y _12948_/C _12950_/Y _12951_/X vssd1 vssd1 vccd1 vccd1 _12955_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11905_ _12018_/A _11905_/B _11905_/C vssd1 vssd1 vccd1 vccd1 _11906_/C sky130_fd_sc_hd__or3_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _15791_/CLK _15673_/D vssd1 vssd1 vccd1 vccd1 _15673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _12885_/A vssd1 vssd1 vccd1 vccd1 _16175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14624_/A _14624_/B _14629_/A vssd1 vssd1 vccd1 vccd1 _16425_/D sky130_fd_sc_hd__nor3_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _16028_/Q _11891_/B _11836_/C vssd1 vssd1 vccd1 vccd1 _11845_/A sky130_fd_sc_hd__and3_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _14555_/A _14555_/B _14555_/C vssd1 vssd1 vccd1 vccd1 _14556_/C sky130_fd_sc_hd__or3_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11776_/A _11767_/B _11767_/C vssd1 vssd1 vccd1 vccd1 _11768_/A sky130_fd_sc_hd__and3_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _16265_/Q _13514_/C _13450_/X vssd1 vssd1 vccd1 vccd1 _13506_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10718_ _10526_/X _10714_/B _10717_/Y vssd1 vssd1 vccd1 vccd1 _15866_/D sky130_fd_sc_hd__o21a_1
X_14486_ _16405_/Q _14486_/B _14486_/C vssd1 vssd1 vccd1 vccd1 _14496_/B sky130_fd_sc_hd__and3_1
X_11698_ _16009_/Q _11922_/B _11698_/C vssd1 vssd1 vccd1 vccd1 _11698_/X sky130_fd_sc_hd__and3_1
X_16225_ _16261_/CLK _16225_/D vssd1 vssd1 vccd1 vccd1 _16225_/Q sky130_fd_sc_hd__dfxtp_1
X_13437_ _13459_/C vssd1 vssd1 vccd1 vccd1 _13473_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10649_ _10649_/A _10649_/B _10649_/C vssd1 vssd1 vccd1 vccd1 _10650_/A sky130_fd_sc_hd__and3_1
XFILLER_127_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16156_ _16555_/Q _16156_/D vssd1 vssd1 vccd1 vccd1 _16156_/Q sky130_fd_sc_hd__dfxtp_1
X_13368_ _13368_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13374_/C sky130_fd_sc_hd__nor2_1
X_15107_ _15180_/A _15107_/B _15111_/B vssd1 vssd1 vccd1 vccd1 _16502_/D sky130_fd_sc_hd__nor3_1
X_12319_ _12320_/B _12320_/C _12320_/A vssd1 vssd1 vccd1 vccd1 _12321_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16087_ _16118_/CLK _16087_/D vssd1 vssd1 vccd1 vccd1 _16087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13299_ _16234_/Q _13467_/B _13305_/C vssd1 vssd1 vccd1 vccd1 _13299_/Y sky130_fd_sc_hd__nand3_1
XFILLER_142_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15038_ _15045_/A _15038_/B _15038_/C vssd1 vssd1 vccd1 vccd1 _15039_/A sky130_fd_sc_hd__and3_1
XFILLER_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07860_ _15588_/Q vssd1 vssd1 vccd1 vccd1 _08295_/A sky130_fd_sc_hd__clkinv_2
XFILLER_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07791_ _07793_/A vssd1 vssd1 vccd1 vccd1 _07791_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16645__50 vssd1 vssd1 vccd1 vccd1 _16645__50/HI _16721_/A sky130_fd_sc_hd__conb_1
XFILLER_84_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09530_ _09750_/A vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _09497_/A _09461_/B _09467_/B vssd1 vssd1 vccd1 vccd1 _15627_/D sky130_fd_sc_hd__nor3_1
XFILLER_64_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08412_ _08430_/A _08430_/B vssd1 vssd1 vccd1 vccd1 _08428_/B sky130_fd_sc_hd__xor2_2
X_09392_ _09301_/X _09390_/B _09304_/X vssd1 vssd1 vccd1 vccd1 _09392_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08343_ _08343_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _08344_/B sky130_fd_sc_hd__xor2_4
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ _08274_/A _08274_/B vssd1 vssd1 vccd1 vccd1 _08275_/B sky130_fd_sc_hd__nor2_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ _16569_/Q _16567_/Q vssd1 vssd1 vccd1 vccd1 _08204_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09728_ _09726_/Y _09733_/A _09722_/C _09723_/C vssd1 vssd1 vccd1 vccd1 _09730_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09659_ _09658_/X _09656_/B _09651_/X vssd1 vssd1 vccd1 vccd1 _09659_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _16145_/Q _12726_/B _12670_/C vssd1 vssd1 vccd1 vccd1 _12670_/Y sky130_fd_sc_hd__nand3_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11737_/A _11621_/B _11621_/C vssd1 vssd1 vccd1 vccd1 _11622_/C sky130_fd_sc_hd__or3_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14340_ _16383_/Q _14380_/C _14339_/X vssd1 vssd1 vccd1 vccd1 _14342_/B sky130_fd_sc_hd__a21oi_1
XFILLER_129_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11552_ _13183_/A vssd1 vssd1 vccd1 vccd1 _15254_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10503_ _15827_/Q _10646_/B _10509_/C vssd1 vssd1 vccd1 vccd1 _10503_/Y sky130_fd_sc_hd__nand3_1
X_11483_ _11491_/A _11483_/B _11483_/C vssd1 vssd1 vccd1 vccd1 _11484_/A sky130_fd_sc_hd__and3_1
X_14271_ _14271_/A _14271_/B vssd1 vssd1 vccd1 vccd1 _14276_/C sky130_fd_sc_hd__nor2_1
X_16010_ _16554_/Q _16010_/D vssd1 vssd1 vccd1 vccd1 _16010_/Q sky130_fd_sc_hd__dfxtp_1
X_13222_ _16224_/Q _13445_/B _13228_/C vssd1 vssd1 vccd1 vccd1 _13224_/C sky130_fd_sc_hd__nand3_1
X_10434_ _15817_/Q _10434_/B _10440_/C vssd1 vssd1 vccd1 vccd1 _10436_/C sky130_fd_sc_hd__nand3_1
XFILLER_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10365_ _10365_/A _10365_/B vssd1 vssd1 vccd1 vccd1 _10366_/B sky130_fd_sc_hd__nor2_1
X_13153_ _13153_/A vssd1 vssd1 vccd1 vccd1 _16213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _12104_/A vssd1 vssd1 vccd1 vccd1 _16065_/D sky130_fd_sc_hd__clkbuf_1
X_13084_ _13084_/A _13084_/B vssd1 vssd1 vccd1 vccd1 _13087_/B sky130_fd_sc_hd__nor2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10290_/C _10291_/C _10293_/Y _10294_/X vssd1 vssd1 vccd1 vccd1 _10297_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_105_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12035_ _12035_/A vssd1 vssd1 vccd1 vccd1 _16055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13986_ _14828_/A vssd1 vssd1 vccd1 vccd1 _13986_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15725_ _15812_/CLK _15725_/D vssd1 vssd1 vccd1 vccd1 _15725_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12937_ _16184_/Q _12945_/C _12879_/X vssd1 vssd1 vccd1 vccd1 _12941_/B sky130_fd_sc_hd__a21o_1
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15656_ _15791_/CLK _15656_/D vssd1 vssd1 vccd1 vccd1 _15656_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _12868_/A _12868_/B _12868_/C vssd1 vssd1 vccd1 vccd1 _12869_/C sky130_fd_sc_hd__or3_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14720_/A _14612_/C vssd1 vssd1 vccd1 vccd1 _14607_/X sky130_fd_sc_hd__or2_1
XFILLER_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11819_ _16026_/Q _11821_/C _11591_/X vssd1 vssd1 vccd1 vccd1 _11819_/Y sky130_fd_sc_hd__a21oi_1
X_15587_ _16551_/CLK _15587_/D vssd1 vssd1 vccd1 vccd1 _15587_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12799_/A _12808_/B vssd1 vssd1 vccd1 vccd1 _12802_/A sky130_fd_sc_hd__or2_1
X_14538_ _16413_/Q _14547_/C _14537_/X vssd1 vssd1 vccd1 vccd1 _14538_/Y sky130_fd_sc_hd__a21oi_1
X_14469_ _14476_/A _14469_/B _14469_/C vssd1 vssd1 vccd1 vccd1 _14470_/A sky130_fd_sc_hd__and3_1
XFILLER_146_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16208_ _16237_/CLK _16208_/D vssd1 vssd1 vccd1 vccd1 _16208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16139_ _16555_/Q _16139_/D vssd1 vssd1 vccd1 vccd1 _16139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08961_ _09294_/A vssd1 vssd1 vccd1 vccd1 _09124_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07912_ _13322_/A _07912_/B vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__xnor2_2
X_08892_ _10285_/C vssd1 vssd1 vccd1 vccd1 _09053_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07843_ input1/X vssd1 vssd1 vccd1 vccd1 _07848_/A sky130_fd_sc_hd__buf_8
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07774_ _07774_/A vssd1 vssd1 vccd1 vccd1 _07774_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09513_ _09513_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09513_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09444_ _15614_/Q _15613_/Q _15612_/Q _09314_/X vssd1 vssd1 vccd1 vccd1 _15624_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _15613_/Q _09382_/C _10750_/B vssd1 vssd1 vccd1 vccd1 _09378_/A sky130_fd_sc_hd__a21oi_1
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08326_ _08326_/A _08137_/A vssd1 vssd1 vccd1 vccd1 _08327_/B sky130_fd_sc_hd__or2b_1
X_08257_ _09220_/C _08076_/B _08075_/A vssd1 vssd1 vccd1 vccd1 _08259_/B sky130_fd_sc_hd__o21a_1
XFILLER_123_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08188_ _08354_/A _08354_/B vssd1 vssd1 vccd1 vccd1 _08189_/B sky130_fd_sc_hd__xnor2_1
XFILLER_146_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ _12968_/A vssd1 vssd1 vccd1 vccd1 _14941_/A sky130_fd_sc_hd__buf_4
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10081_ _10081_/A _10081_/B _10081_/C vssd1 vssd1 vccd1 vccd1 _10082_/C sky130_fd_sc_hd__nand3_1
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13840_ _13927_/A _13840_/B _13844_/A vssd1 vssd1 vccd1 vccd1 _16310_/D sky130_fd_sc_hd__nor3_1
XFILLER_75_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13771_ _13881_/A vssd1 vssd1 vccd1 vccd1 _13811_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10983_ _11266_/A vssd1 vssd1 vccd1 vccd1 _11097_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15510_ _16551_/CLK _15510_/D vssd1 vssd1 vccd1 vccd1 _15510_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12722_ _12722_/A vssd1 vssd1 vccd1 vccd1 _16152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16490_ _16607_/CLK _16490_/D vssd1 vssd1 vccd1 vccd1 _16490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15441_ _16357_/Q _16356_/Q _16355_/Q _15440_/X vssd1 vssd1 vccd1 vccd1 _16615_/D
+ sky130_fd_sc_hd__o31a_1
X_12653_ _12653_/A _12653_/B _12659_/A vssd1 vssd1 vccd1 vccd1 _16142_/D sky130_fd_sc_hd__nor3_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _11604_/A _11604_/B _11604_/C vssd1 vssd1 vccd1 vccd1 _11605_/A sky130_fd_sc_hd__and3_1
X_15372_ _15378_/A vssd1 vssd1 vccd1 vccd1 _15372_/X sky130_fd_sc_hd__buf_2
X_12584_ _12751_/A vssd1 vssd1 vccd1 vccd1 _12625_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14323_ _16381_/Q _14486_/B _14323_/C vssd1 vssd1 vccd1 vccd1 _14332_/B sky130_fd_sc_hd__and3_1
X_11535_ _15986_/Q _11644_/B _11536_/C vssd1 vssd1 vccd1 vccd1 _11535_/X sky130_fd_sc_hd__and3_1
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14254_ _14250_/Y _14252_/X _14253_/Y _14248_/C vssd1 vssd1 vccd1 vccd1 _14256_/B
+ sky130_fd_sc_hd__o211ai_1
X_11466_ _11467_/B _11467_/C _11467_/A vssd1 vssd1 vccd1 vccd1 _11468_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ _13317_/A vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10417_ _10220_/X _10409_/B _10412_/B _10416_/Y vssd1 vssd1 vccd1 vccd1 _15811_/D
+ sky130_fd_sc_hd__o31a_1
X_11397_ _16567_/Q vssd1 vssd1 vccd1 vccd1 _11412_/C sky130_fd_sc_hd__inv_2
X_14185_ _16362_/Q _14185_/B _14187_/C vssd1 vssd1 vccd1 vccd1 _14185_/X sky130_fd_sc_hd__and3_1
XFILLER_99_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13136_ _16211_/Q _13194_/B _13143_/C vssd1 vssd1 vccd1 vccd1 _13136_/Y sky130_fd_sc_hd__nand3_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _15801_/Q _10446_/B _10355_/C vssd1 vssd1 vccd1 vccd1 _10348_/X sky130_fd_sc_hd__and3_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _15776_/Q _15775_/Q _15774_/Q _10227_/X vssd1 vssd1 vccd1 vccd1 _15786_/D
+ sky130_fd_sc_hd__o31a_1
X_13067_ _16203_/Q _13076_/C _12901_/X vssd1 vssd1 vccd1 vccd1 _13067_/Y sky130_fd_sc_hd__a21oi_1
X_12018_ _12018_/A _12018_/B _12018_/C vssd1 vssd1 vccd1 vccd1 _12019_/C sky130_fd_sc_hd__or3_1
XFILLER_120_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16757_ _16757_/A _07776_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
X_13969_ _13977_/A _13969_/B _13969_/C vssd1 vssd1 vccd1 vccd1 _13970_/A sky130_fd_sc_hd__and3_1
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15708_ _15812_/CLK _15708_/D vssd1 vssd1 vccd1 vccd1 _15708_/Q sky130_fd_sc_hd__dfxtp_2
X_16688_ _16688_/A _07785_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _15791_/CLK _15639_/D vssd1 vssd1 vccd1 vccd1 _15639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09160_ _09240_/A _09165_/C vssd1 vssd1 vccd1 vccd1 _09162_/A sky130_fd_sc_hd__and2_1
X_08111_ _08766_/C _08111_/B vssd1 vssd1 vccd1 vccd1 _08111_/X sky130_fd_sc_hd__or2_1
XFILLER_147_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09091_ _15542_/Q _15541_/Q _15540_/Q _09090_/X vssd1 vssd1 vccd1 vccd1 _15552_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ _16451_/Q vssd1 vssd1 vccd1 vccd1 _14675_/A sky130_fd_sc_hd__inv_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09993_ _09994_/B _09994_/C _09994_/A vssd1 vssd1 vccd1 vccd1 _09995_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08944_ _08942_/Y _08950_/A _08939_/C _08940_/C vssd1 vssd1 vccd1 vccd1 _08946_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08875_ _08872_/X _08867_/B _08870_/B _08874_/Y vssd1 vssd1 vccd1 vccd1 _15503_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07826_ _07830_/A vssd1 vssd1 vccd1 vccd1 _07826_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07757_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07762_/A sky130_fd_sc_hd__buf_12
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ _09423_/A _09422_/Y _09423_/B vssd1 vssd1 vccd1 vccd1 _09427_/Y sky130_fd_sc_hd__o21bai_1
X_09358_ _09371_/C vssd1 vssd1 vccd1 vccd1 _09382_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08309_ _15293_/C _08309_/B vssd1 vssd1 vccd1 vccd1 _08309_/Y sky130_fd_sc_hd__xnor2_1
X_09289_ _09282_/Y _09288_/X _09129_/X vssd1 vssd1 vccd1 vccd1 _09289_/Y sky130_fd_sc_hd__a21oi_1
X_11320_ _11320_/A vssd1 vssd1 vccd1 vccd1 _15954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11251_ _15946_/Q _11253_/C _11023_/X vssd1 vssd1 vccd1 vccd1 _11251_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10202_ _10202_/A vssd1 vssd1 vccd1 vccd1 _15772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11182_ _15936_/Q _11190_/C _11181_/X vssd1 vssd1 vccd1 vccd1 _11185_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10133_ _15764_/Q _10190_/B _10133_/C vssd1 vssd1 vccd1 vccd1 _10133_/X sky130_fd_sc_hd__and3_1
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15990_ _16005_/CLK _15990_/D vssd1 vssd1 vccd1 vccd1 _15990_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_85_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10064_ _10058_/B _10062_/B _09125_/A vssd1 vssd1 vccd1 vccd1 _10065_/B sky130_fd_sc_hd__o21a_1
X_14941_ _14941_/A vssd1 vssd1 vccd1 vccd1 _15156_/B sky130_fd_sc_hd__buf_2
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14872_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14872_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16611_ input11/X _16611_/D vssd1 vssd1 vccd1 vccd1 _16611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13823_ _13823_/A _13831_/B vssd1 vssd1 vccd1 vccd1 _13825_/A sky130_fd_sc_hd__or2_1
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16542_ _16595_/CLK _16542_/D vssd1 vssd1 vccd1 vccd1 _16711_/A sky130_fd_sc_hd__dfxtp_4
X_13754_ _13751_/Y _13752_/X _13753_/Y _13748_/C vssd1 vssd1 vccd1 vccd1 _13756_/B
+ sky130_fd_sc_hd__o211ai_1
X_10966_ _10981_/A _10966_/B _10966_/C vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__and3_1
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _12718_/C vssd1 vssd1 vccd1 vccd1 _12726_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16473_ _16607_/CLK _16473_/D vssd1 vssd1 vccd1 vccd1 _16473_/Q sky130_fd_sc_hd__dfxtp_1
X_13685_ _13681_/Y _13683_/X _13684_/Y _13679_/C vssd1 vssd1 vccd1 vccd1 _13687_/B
+ sky130_fd_sc_hd__o211ai_1
X_10897_ _12655_/A vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__clkbuf_4
X_15424_ _16245_/Q _16244_/Q _16243_/Q _15422_/X vssd1 vssd1 vccd1 vccd1 _16601_/D
+ sky130_fd_sc_hd__o31a_1
X_12636_ _12636_/A _12636_/B vssd1 vssd1 vccd1 vccd1 _12637_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15355_ _15355_/A _15358_/C vssd1 vssd1 vccd1 vccd1 _15357_/A sky130_fd_sc_hd__and2_1
X_12567_ _12567_/A vssd1 vssd1 vccd1 vccd1 _12567_/X sky130_fd_sc_hd__buf_2
X_14306_ _14314_/A _14306_/B _14306_/C vssd1 vssd1 vccd1 vccd1 _14307_/A sky130_fd_sc_hd__and3_1
X_11518_ _15983_/Q _11560_/C _11517_/X vssd1 vssd1 vccd1 vccd1 _11520_/B sky130_fd_sc_hd__a21oi_1
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15286_ _15293_/C _15286_/B vssd1 vssd1 vccd1 vccd1 _15286_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_144_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _12505_/A _12498_/B _12498_/C vssd1 vssd1 vccd1 vccd1 _12499_/A sky130_fd_sc_hd__and3_1
X_14237_ _16369_/Q _14458_/B _14237_/C vssd1 vssd1 vccd1 vccd1 _14237_/X sky130_fd_sc_hd__and3_1
X_11449_ _11447_/A _11447_/B _11448_/X vssd1 vssd1 vccd1 vccd1 _15972_/D sky130_fd_sc_hd__a21oi_1
XFILLER_125_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14168_ _14201_/C vssd1 vssd1 vccd1 vccd1 _14207_/C sky130_fd_sc_hd__clkbuf_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _16210_/Q _13342_/B _13120_/C vssd1 vssd1 vccd1 vccd1 _13119_/X sky130_fd_sc_hd__and3_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14099_ _14205_/A _14099_/B _14103_/B vssd1 vssd1 vccd1 vccd1 _16347_/D sky130_fd_sc_hd__nor3_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08660_ _09792_/A vssd1 vssd1 vccd1 vccd1 _10276_/A sky130_fd_sc_hd__buf_4
XFILLER_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08591_ _08592_/B _08592_/C _08592_/A vssd1 vssd1 vccd1 vccd1 _08593_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09212_ _15584_/Q _09231_/C _09051_/X vssd1 vssd1 vccd1 vccd1 _09214_/B sky130_fd_sc_hd__a21oi_1
XFILLER_61_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09143_ _09143_/A vssd1 vssd1 vccd1 vccd1 _15563_/D sky130_fd_sc_hd__clkbuf_1
X_09074_ _09074_/A _09074_/B vssd1 vssd1 vccd1 vccd1 _09074_/X sky130_fd_sc_hd__or2_1
XFILLER_107_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08025_ _15849_/Q _15831_/Q vssd1 vssd1 vccd1 vccd1 _08217_/A sky130_fd_sc_hd__nand2_1
XFILLER_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09976_ _09749_/X _09973_/B _09975_/Y vssd1 vssd1 vccd1 vccd1 _15730_/D sky130_fd_sc_hd__o21a_1
XFILLER_77_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08927_ _15350_/A vssd1 vssd1 vccd1 vccd1 _08927_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08858_ _10492_/A vssd1 vssd1 vccd1 vccd1 _10447_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07809_ _07811_/A vssd1 vssd1 vccd1 vccd1 _07809_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08789_ _08644_/X _08791_/C _08708_/X vssd1 vssd1 vccd1 vccd1 _08790_/B sky130_fd_sc_hd__o21ai_1
XFILLER_72_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10820_ _11957_/A vssd1 vssd1 vccd1 vccd1 _11051_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10751_ _10748_/Y _10757_/A _10750_/Y _10746_/C vssd1 vssd1 vccd1 vccd1 _10753_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _13470_/A _13470_/B _13470_/C vssd1 vssd1 vccd1 vccd1 _13471_/A sky130_fd_sc_hd__and3_1
XFILLER_139_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ _10738_/A _10682_/B _10682_/C vssd1 vssd1 vccd1 vccd1 _10683_/A sky130_fd_sc_hd__and3_1
X_12421_ _16585_/Q vssd1 vssd1 vccd1 vccd1 _12435_/C sky130_fd_sc_hd__inv_2
XFILLER_139_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15140_ _16510_/Q _15142_/C _14979_/X vssd1 vssd1 vccd1 vccd1 _15140_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12352_ _16101_/Q _12516_/B _12352_/C vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__and3_1
XFILLER_5_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11303_ _11297_/C _11298_/C _11300_/Y _11301_/X vssd1 vssd1 vccd1 vccd1 _11304_/C
+ sky130_fd_sc_hd__a211o_1
X_15071_ _15090_/C vssd1 vssd1 vccd1 vccd1 _15103_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12283_ _12283_/A _12283_/B _12283_/C vssd1 vssd1 vccd1 vccd1 _12284_/A sky130_fd_sc_hd__and3_1
X_14022_ _16338_/Q _14024_/C _13853_/X vssd1 vssd1 vccd1 vccd1 _14022_/Y sky130_fd_sc_hd__a21oi_1
X_11234_ _15943_/Q _11275_/C _11233_/X vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__a21oi_1
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11165_ _11332_/A _11169_/C vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__or2_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10116_ _09207_/X _10114_/B _10012_/X vssd1 vssd1 vccd1 vccd1 _10116_/Y sky130_fd_sc_hd__a21oi_1
X_15973_ _16005_/CLK _15973_/D vssd1 vssd1 vccd1 vccd1 _15973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11096_ _11094_/Y _11088_/C _11090_/Y _11101_/A vssd1 vssd1 vccd1 vccd1 _11101_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_103_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10047_ _10045_/Y _10041_/C _10043_/Y _10044_/X vssd1 vssd1 vccd1 vccd1 _10048_/C
+ sky130_fd_sc_hd__a211o_1
X_14924_ _16474_/Q _15033_/B _14925_/C vssd1 vssd1 vccd1 vccd1 _14924_/X sky130_fd_sc_hd__and3_1
XFILLER_76_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14855_ _14855_/A _14855_/B _14855_/C vssd1 vssd1 vccd1 vccd1 _14856_/C sky130_fd_sc_hd__nand3_1
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13806_ _16307_/Q _13914_/B _13815_/C vssd1 vssd1 vccd1 vccd1 _13806_/X sky130_fd_sc_hd__and3_1
XFILLER_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14786_ _14800_/C vssd1 vssd1 vccd1 vccd1 _14808_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11998_ _11998_/A _11998_/B _11998_/C vssd1 vssd1 vccd1 vccd1 _11999_/A sky130_fd_sc_hd__and3_1
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16525_ _16595_/CLK _16525_/D vssd1 vssd1 vccd1 vccd1 _16525_/Q sky130_fd_sc_hd__dfxtp_1
X_13737_ _16297_/Q _13745_/C _13736_/X vssd1 vssd1 vccd1 vccd1 _13737_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10949_ _10970_/C vssd1 vssd1 vccd1 vccd1 _10985_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16456_ _16607_/CLK _16456_/D vssd1 vssd1 vccd1 vccd1 _16456_/Q sky130_fd_sc_hd__dfxtp_1
X_13668_ _16288_/Q _13731_/B _13676_/C vssd1 vssd1 vccd1 vccd1 _13670_/C sky130_fd_sc_hd__nand3_1
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15407_ _16141_/Q _16140_/Q _16139_/Q _15403_/X vssd1 vssd1 vccd1 vccd1 _16588_/D
+ sky130_fd_sc_hd__o31a_1
X_12619_ _12901_/A vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__buf_2
X_16387_ _16389_/CLK _16387_/D vssd1 vssd1 vccd1 vccd1 _16387_/Q sky130_fd_sc_hd__dfxtp_1
X_13599_ _13600_/B _13600_/C _13546_/X vssd1 vssd1 vccd1 vccd1 _13601_/B sky130_fd_sc_hd__o21ai_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15338_ _15338_/A _15338_/B _15338_/C vssd1 vssd1 vccd1 vccd1 _15339_/A sky130_fd_sc_hd__and3_1
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_0 _07805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15269_ _15269_/A _15269_/B vssd1 vssd1 vccd1 vccd1 _15270_/B sky130_fd_sc_hd__nor2_1
XFILLER_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09830_ _09828_/Y _09819_/C _09822_/Y _09826_/X vssd1 vssd1 vccd1 vccd1 _09831_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _15691_/Q _09945_/B _09761_/C vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__and3_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08712_ _08663_/X _08710_/A _08711_/X vssd1 vssd1 vccd1 vccd1 _08712_/Y sky130_fd_sc_hd__a21oi_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _15677_/Q _09692_/B _09692_/C vssd1 vssd1 vccd1 vccd1 _09692_/X sky130_fd_sc_hd__and3_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08643_ _10016_/A vssd1 vssd1 vccd1 vccd1 _09038_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _12932_/A vssd1 vssd1 vccd1 vccd1 _14906_/A sky130_fd_sc_hd__buf_6
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ _09126_/A vssd1 vssd1 vccd1 vccd1 _09126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09057_ _15549_/Q _09220_/B _09057_/C vssd1 vssd1 vccd1 vccd1 _09059_/C sky130_fd_sc_hd__nand3_1
XFILLER_2_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08008_ _16617_/Q vssd1 vssd1 vccd1 vccd1 _14222_/A sky130_fd_sc_hd__inv_4
XFILLER_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09959_ _15730_/Q _09966_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _09962_/A sky130_fd_sc_hd__a21oi_1
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12970_ _16187_/Q _13194_/B _12975_/C vssd1 vssd1 vccd1 vccd1 _12970_/Y sky130_fd_sc_hd__nand3_1
XFILLER_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11921_ _16041_/Q _11930_/C _11755_/X vssd1 vssd1 vccd1 vccd1 _11921_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14640_ _16428_/Q _14697_/B _14640_/C vssd1 vssd1 vccd1 vccd1 _14640_/Y sky130_fd_sc_hd__nand3_1
XFILLER_122_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11852_ _12018_/A _11852_/B _11852_/C vssd1 vssd1 vccd1 vccd1 _11853_/C sky130_fd_sc_hd__or3_1
XFILLER_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10803_ _15883_/Q _10812_/C _10755_/B vssd1 vssd1 vccd1 vccd1 _10803_/Y sky130_fd_sc_hd__a21oi_1
X_14571_ _14571_/A _14571_/B _14571_/C vssd1 vssd1 vccd1 vccd1 _14572_/C sky130_fd_sc_hd__nand3_1
X_11783_ _11805_/A _11783_/B _11787_/B vssd1 vssd1 vccd1 vccd1 _16019_/D sky130_fd_sc_hd__nor3_1
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16310_ _16346_/CLK _16310_/D vssd1 vssd1 vccd1 vccd1 _16310_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13522_ _14647_/A vssd1 vssd1 vccd1 vccd1 _13753_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10734_ _15872_/Q _10735_/C _09416_/B vssd1 vssd1 vccd1 vccd1 _10734_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_14_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16241_ _16261_/CLK _16241_/D vssd1 vssd1 vccd1 vccd1 _16241_/Q sky130_fd_sc_hd__dfxtp_1
X_13453_ _13451_/Y _13452_/X _13447_/C _13448_/C vssd1 vssd1 vccd1 vccd1 _13455_/B
+ sky130_fd_sc_hd__o211ai_1
X_10665_ _15353_/A _10665_/B vssd1 vssd1 vccd1 vccd1 _10665_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ _16107_/Q _12629_/B _12409_/C vssd1 vssd1 vccd1 vccd1 _12404_/Y sky130_fd_sc_hd__nand3_1
X_16172_ _16555_/Q _16172_/D vssd1 vssd1 vccd1 vccd1 _16172_/Q sky130_fd_sc_hd__dfxtp_1
X_13384_ _13498_/A _13384_/B _13388_/A vssd1 vssd1 vccd1 vccd1 _16246_/D sky130_fd_sc_hd__nor3_1
X_10596_ _10649_/A _10596_/B _10596_/C vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__and3_1
XFILLER_139_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15123_ _15142_/C vssd1 vssd1 vccd1 vccd1 _15155_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12335_ _12343_/A _12335_/B _12335_/C vssd1 vssd1 vccd1 vccd1 _12336_/A sky130_fd_sc_hd__and3_1
XFILLER_127_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15054_ _16495_/Q _15055_/C _14828_/X vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__a21oi_1
XFILLER_99_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12266_ _12283_/A _12266_/B _12266_/C vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__and3_1
XFILLER_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14005_ _14848_/A vssd1 vssd1 vccd1 vccd1 _14227_/B sky130_fd_sc_hd__clkbuf_2
X_11217_ _15941_/Q _11381_/B _11217_/C vssd1 vssd1 vccd1 vccd1 _11226_/B sky130_fd_sc_hd__and3_1
X_12197_ _16080_/Q _12204_/C _12029_/X vssd1 vssd1 vccd1 vccd1 _12200_/B sky130_fd_sc_hd__a21o_1
X_11148_ _11148_/A _11148_/B _11148_/C vssd1 vssd1 vccd1 vccd1 _11149_/A sky130_fd_sc_hd__and3_1
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15956_ _16005_/CLK _15956_/D vssd1 vssd1 vccd1 vccd1 _15956_/Q sky130_fd_sc_hd__dfxtp_1
X_11079_ _11075_/Y _11076_/X _11078_/Y _11073_/C vssd1 vssd1 vccd1 vccd1 _11081_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_110_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14907_ _16471_/Q _14947_/C _14906_/X vssd1 vssd1 vccd1 vccd1 _14909_/B sky130_fd_sc_hd__a21oi_1
X_15887_ _16553_/Q _15887_/D vssd1 vssd1 vccd1 vccd1 _15887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14838_ _14839_/B _14839_/C _14669_/X vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__o21ai_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14769_ _16450_/Q _14770_/C _14544_/X vssd1 vssd1 vccd1 vccd1 _14771_/A sky130_fd_sc_hd__a21oi_1
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ _16607_/CLK _16508_/D vssd1 vssd1 vccd1 vccd1 _16508_/Q sky130_fd_sc_hd__dfxtp_1
X_08290_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08291_/B sky130_fd_sc_hd__xor2_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16439_ _16595_/CLK _16439_/D vssd1 vssd1 vccd1 vccd1 _16439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09813_ _10492_/A vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__buf_2
XFILLER_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09744_ _09744_/A vssd1 vssd1 vccd1 vccd1 _09744_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09675_ _09810_/A _09675_/B _09675_/C vssd1 vssd1 vccd1 vccd1 _09676_/A sky130_fd_sc_hd__and3_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _14872_/A vssd1 vssd1 vccd1 vccd1 _10456_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _08545_/A _08545_/B _08556_/X vssd1 vssd1 vccd1 vccd1 _08567_/A sky130_fd_sc_hd__a21oi_2
XFILLER_23_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08488_ _15304_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08489_/A sky130_fd_sc_hd__and2_1
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10450_ _10448_/Y _10443_/C _10445_/Y _10446_/X vssd1 vssd1 vccd1 vccd1 _10451_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09109_ _15560_/Q _09110_/C _08989_/X vssd1 vssd1 vccd1 vccd1 _09111_/A sky130_fd_sc_hd__a21oi_1
X_10381_ _15808_/Q _10388_/C _10181_/X vssd1 vssd1 vccd1 vccd1 _10384_/B sky130_fd_sc_hd__a21o_1
X_12120_ _16067_/Q _12347_/B _12125_/C vssd1 vssd1 vccd1 vccd1 _12120_/Y sky130_fd_sc_hd__nand3_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12051_ _16059_/Q _12059_/C _12050_/X vssd1 vssd1 vccd1 vccd1 _12051_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ _11036_/A _11002_/B _11002_/C vssd1 vssd1 vccd1 vccd1 _11003_/A sky130_fd_sc_hd__and3_1
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15810_ _15812_/CLK _15810_/D vssd1 vssd1 vccd1 vccd1 _15810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15741_ _16551_/CLK _15741_/D vssd1 vssd1 vccd1 vccd1 _15741_/Q sky130_fd_sc_hd__dfxtp_1
X_12953_ _12950_/Y _12951_/X _12952_/Y _12948_/C vssd1 vssd1 vccd1 vccd1 _12955_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11904_ _11905_/B _11905_/C _11850_/X vssd1 vssd1 vccd1 vccd1 _11906_/B sky130_fd_sc_hd__o21ai_1
X_15672_ _15791_/CLK _15672_/D vssd1 vssd1 vccd1 vccd1 _15672_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12907_/A _12884_/B _12884_/C vssd1 vssd1 vccd1 vccd1 _12885_/A sky130_fd_sc_hd__and3_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14623_ _16426_/Q _14790_/B _14633_/C vssd1 vssd1 vccd1 vccd1 _14629_/A sky130_fd_sc_hd__and3_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _16028_/Q _11843_/C _11719_/X vssd1 vssd1 vccd1 vccd1 _11835_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14555_/B _14555_/C _14387_/X vssd1 vssd1 vccd1 vccd1 _14556_/B sky130_fd_sc_hd__o21ai_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11764_/Y _11760_/C _11762_/Y _11763_/X vssd1 vssd1 vccd1 vccd1 _11767_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13505_/A vssd1 vssd1 vccd1 vccd1 _16263_/D sky130_fd_sc_hd__clkbuf_1
X_10717_ _09308_/X _10714_/B _10716_/X vssd1 vssd1 vccd1 vccd1 _10717_/Y sky130_fd_sc_hd__a21oi_1
X_14485_ _16405_/Q _14486_/C _14265_/X vssd1 vssd1 vccd1 vccd1 _14487_/A sky130_fd_sc_hd__a21oi_1
X_11697_ _11978_/A vssd1 vssd1 vccd1 vccd1 _11922_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16224_ _16261_/CLK _16224_/D vssd1 vssd1 vccd1 vccd1 _16224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13436_ _13452_/C vssd1 vssd1 vccd1 vccd1 _13459_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10648_ _10646_/Y _10642_/C _10644_/Y _10645_/X vssd1 vssd1 vccd1 vccd1 _10649_/C
+ sky130_fd_sc_hd__a211o_1
X_16155_ _16555_/Q _16155_/D vssd1 vssd1 vccd1 vccd1 _16155_/Q sky130_fd_sc_hd__dfxtp_1
X_13367_ _14210_/A vssd1 vssd1 vccd1 vccd1 _13596_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10579_ _10583_/C vssd1 vssd1 vccd1 vccd1 _10593_/C sky130_fd_sc_hd__clkbuf_1
X_15106_ _15104_/Y _15100_/C _15102_/Y _15111_/A vssd1 vssd1 vccd1 vccd1 _15111_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_142_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ _16096_/Q _12318_/B _12325_/C vssd1 vssd1 vccd1 vccd1 _12320_/C sky130_fd_sc_hd__nand3_1
X_16086_ _16118_/CLK _16086_/D vssd1 vssd1 vccd1 vccd1 _16086_/Q sky130_fd_sc_hd__dfxtp_2
X_13298_ _16235_/Q _13350_/B _13305_/C vssd1 vssd1 vccd1 vccd1 _13298_/X sky130_fd_sc_hd__and3_1
X_15037_ _15035_/Y _15030_/C _15032_/Y _15033_/X vssd1 vssd1 vccd1 vccd1 _15038_/C
+ sky130_fd_sc_hd__a211o_1
X_12249_ _12271_/C vssd1 vssd1 vccd1 vccd1 _12287_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07790_ _07793_/A vssd1 vssd1 vccd1 vccd1 _07790_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15939_ _15365_/A _15939_/D vssd1 vssd1 vccd1 vccd1 _15939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09460_ _09453_/C _09454_/C _09456_/Y _09467_/A vssd1 vssd1 vccd1 vccd1 _09467_/B
+ sky130_fd_sc_hd__a211oi_1
X_16660__65 vssd1 vssd1 vccd1 vccd1 _16660__65/HI _16736_/A sky130_fd_sc_hd__conb_1
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08411_ _08411_/A _08431_/A vssd1 vssd1 vccd1 vccd1 _08430_/B sky130_fd_sc_hd__xnor2_2
X_09391_ _09291_/X _09389_/B _09390_/Y vssd1 vssd1 vccd1 vccd1 _15612_/D sky130_fd_sc_hd__o21a_1
XFILLER_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08342_ _08435_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__xor2_4
XFILLER_149_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08273_ _08273_/A _08273_/B vssd1 vssd1 vccd1 vccd1 _08274_/B sky130_fd_sc_hd__and2_1
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07988_ _16569_/Q _16567_/Q vssd1 vssd1 vccd1 vccd1 _07991_/B sky130_fd_sc_hd__or2_1
XFILLER_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09727_ _15684_/Q _09914_/B _09727_/C vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__and3_1
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09658_ _10469_/A vssd1 vssd1 vccd1 vccd1 _09658_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08609_ _08605_/Y _08621_/A _08592_/C _08593_/C vssd1 vssd1 vccd1 vccd1 _08611_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09589_/A vssd1 vssd1 vccd1 vccd1 _15653_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11621_/B _11621_/C _11567_/X vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__o21ai_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11551_ _15988_/Q _11607_/B _11551_/C vssd1 vssd1 vccd1 vccd1 _11562_/A sky130_fd_sc_hd__and3_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10502_ _15828_/Q _10691_/B _10509_/C vssd1 vssd1 vccd1 vccd1 _10502_/X sky130_fd_sc_hd__and3_1
X_14270_ _14270_/A _14270_/B vssd1 vssd1 vccd1 vccd1 _14271_/B sky130_fd_sc_hd__nor2_1
X_11482_ _11480_/Y _11476_/C _11478_/Y _11479_/X vssd1 vssd1 vccd1 vccd1 _11483_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13221_ _13786_/A vssd1 vssd1 vccd1 vccd1 _13445_/B sky130_fd_sc_hd__clkbuf_2
X_10433_ _15817_/Q _10440_/C _10432_/X vssd1 vssd1 vccd1 vccd1 _10436_/B sky130_fd_sc_hd__a21o_1
XFILLER_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13152_ _13190_/A _13152_/B _13152_/C vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__and3_1
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10364_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10365_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _12113_/A _12103_/B _12103_/C vssd1 vssd1 vccd1 vccd1 _12104_/A sky130_fd_sc_hd__and3_1
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13083_/A _13093_/B vssd1 vssd1 vccd1 vccd1 _13087_/A sky130_fd_sc_hd__or2_1
X_10295_ _10293_/Y _10294_/X _10290_/C _10291_/C vssd1 vssd1 vccd1 vccd1 _10297_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_3_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12034_ _12056_/A _12034_/B _12034_/C vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__and3_1
XFILLER_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13985_ _14063_/A _13985_/B _13991_/B vssd1 vssd1 vccd1 vccd1 _16331_/D sky130_fd_sc_hd__nor3_1
XFILLER_19_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15724_ _15812_/CLK _15724_/D vssd1 vssd1 vccd1 vccd1 _15724_/Q sky130_fd_sc_hd__dfxtp_2
X_12936_ _12936_/A _12936_/B _12941_/A vssd1 vssd1 vccd1 vccd1 _16182_/D sky130_fd_sc_hd__nor3_1
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15655_ _15791_/CLK _15655_/D vssd1 vssd1 vccd1 vccd1 _15655_/Q sky130_fd_sc_hd__dfxtp_1
X_12867_ _12868_/B _12868_/C _12699_/X vssd1 vssd1 vccd1 vccd1 _12869_/B sky130_fd_sc_hd__o21ai_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _11818_/A vssd1 vssd1 vccd1 vccd1 _16024_/D sky130_fd_sc_hd__clkbuf_1
X_14606_ _14606_/A _14606_/B vssd1 vssd1 vccd1 vccd1 _14612_/C sky130_fd_sc_hd__nor2_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15586_ _16551_/CLK _15586_/D vssd1 vssd1 vccd1 vccd1 _15586_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _16165_/Q _12798_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12808_/B sky130_fd_sc_hd__and3_1
XFILLER_14_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14537_/X sky130_fd_sc_hd__buf_2
X_11749_ _16016_/Q _11757_/C _11748_/X vssd1 vssd1 vccd1 vccd1 _11752_/B sky130_fd_sc_hd__a21o_1
X_14468_ _14466_/Y _14461_/C _14463_/Y _14464_/X vssd1 vssd1 vccd1 vccd1 _14469_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_146_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16207_ _16237_/CLK _16207_/D vssd1 vssd1 vccd1 vccd1 _16207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13419_ _13417_/Y _13412_/C _13415_/Y _13426_/A vssd1 vssd1 vccd1 vccd1 _13426_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_127_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14399_ _16392_/Q _14406_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14402_/B sky130_fd_sc_hd__a21o_1
X_16138_ _16555_/Q _16138_/D vssd1 vssd1 vccd1 vccd1 _16138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08960_ _08960_/A _08960_/B vssd1 vssd1 vccd1 vccd1 _15522_/D sky130_fd_sc_hd__nor2_1
X_16069_ _16554_/Q _16069_/D vssd1 vssd1 vccd1 vccd1 _16069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07911_ _13943_/A _07911_/B vssd1 vssd1 vccd1 vccd1 _07912_/B sky130_fd_sc_hd__xnor2_4
X_08891_ _15512_/Q _08907_/C _08843_/X vssd1 vssd1 vccd1 vccd1 _08894_/B sky130_fd_sc_hd__a21oi_1
XFILLER_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07842_ _07842_/A vssd1 vssd1 vccd1 vccd1 _07842_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07773_ _07774_/A vssd1 vssd1 vccd1 vccd1 _07773_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09512_ _15640_/Q _09641_/B _09519_/C vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__and3_1
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _09443_/A _09443_/B vssd1 vssd1 vccd1 vccd1 _15623_/D sky130_fd_sc_hd__nor2_1
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ _09374_/A _09374_/B _09377_/B vssd1 vssd1 vccd1 vccd1 _15609_/D sky130_fd_sc_hd__nor3_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08325_ _08325_/A _08136_/A vssd1 vssd1 vccd1 vccd1 _08327_/A sky130_fd_sc_hd__or2b_1
X_08256_ _08256_/A vssd1 vssd1 vccd1 vccd1 _09220_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_08187_ _08355_/A _08187_/B vssd1 vssd1 vccd1 vccd1 _08354_/B sky130_fd_sc_hd__and2_1
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10080_ _10081_/B _10081_/C _10081_/A vssd1 vssd1 vccd1 vccd1 _10082_/B sky130_fd_sc_hd__a21o_1
XFILLER_102_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13770_ _13768_/A _13768_/B _13769_/X vssd1 vssd1 vccd1 vccd1 _16300_/D sky130_fd_sc_hd__a21oi_1
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10982_ _10982_/A vssd1 vssd1 vccd1 vccd1 _15906_/D sky130_fd_sc_hd__clkbuf_1
X_12721_ _12736_/A _12721_/B _12721_/C vssd1 vssd1 vccd1 vccd1 _12722_/A sky130_fd_sc_hd__and3_1
XFILLER_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15440_ _15440_/A vssd1 vssd1 vccd1 vccd1 _15440_/X sky130_fd_sc_hd__clkbuf_2
X_12652_ _16143_/Q _12818_/B _12663_/C vssd1 vssd1 vccd1 vccd1 _12659_/A sky130_fd_sc_hd__and3_1
XFILLER_31_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _11601_/Y _11597_/C _11599_/Y _11600_/X vssd1 vssd1 vccd1 vccd1 _11604_/C
+ sky130_fd_sc_hd__a211o_1
X_15371_ _15909_/Q _15908_/Q _15907_/Q _15363_/X vssd1 vssd1 vccd1 vccd1 _16559_/D
+ sky130_fd_sc_hd__o31a_1
X_12583_ _12581_/A _12581_/B _12582_/X vssd1 vssd1 vccd1 vccd1 _16132_/D sky130_fd_sc_hd__a21oi_1
X_14322_ _16381_/Q _14323_/C _14265_/X vssd1 vssd1 vccd1 vccd1 _14324_/A sky130_fd_sc_hd__a21oi_1
X_11534_ _15986_/Q _11536_/C _11306_/X vssd1 vssd1 vccd1 vccd1 _11534_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14253_ _16370_/Q _14311_/B _14260_/C vssd1 vssd1 vccd1 vccd1 _14253_/Y sky130_fd_sc_hd__nand3_1
X_11465_ _15976_/Q _11465_/B _11473_/C vssd1 vssd1 vccd1 vccd1 _11467_/C sky130_fd_sc_hd__nand3_1
XFILLER_125_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _13202_/A _13202_/B _13203_/X vssd1 vssd1 vccd1 vccd1 _16220_/D sky130_fd_sc_hd__a21oi_1
X_10416_ _10573_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10416_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14184_ _16362_/Q _14187_/C _14132_/X vssd1 vssd1 vccd1 vccd1 _14184_/Y sky130_fd_sc_hd__a21oi_1
X_11396_ _11963_/A vssd1 vssd1 vccd1 vccd1 _11520_/A sky130_fd_sc_hd__buf_2
X_13135_ _16212_/Q _13305_/B _13135_/C vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__and3_1
X_10347_ _15801_/Q _10355_/C _10138_/X vssd1 vssd1 vccd1 vccd1 _10347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13066_ _13066_/A vssd1 vssd1 vccd1 vccd1 _16201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10278_ _10276_/X _10274_/B _10277_/Y vssd1 vssd1 vccd1 vccd1 _15785_/D sky130_fd_sc_hd__o21a_1
XFILLER_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12017_ _12018_/B _12018_/C _11850_/X vssd1 vssd1 vccd1 vccd1 _12019_/B sky130_fd_sc_hd__o21ai_1
XFILLER_66_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16756_ _16756_/A _07774_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
X_13968_ _13966_/Y _13961_/C _13963_/Y _13965_/X vssd1 vssd1 vccd1 vccd1 _13969_/C
+ sky130_fd_sc_hd__a211o_1
X_15707_ _15812_/CLK _15707_/D vssd1 vssd1 vccd1 vccd1 _15707_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12919_ _12919_/A _12919_/B vssd1 vssd1 vccd1 vccd1 _12925_/C sky130_fd_sc_hd__nor2_1
X_13899_ _16321_/Q _13908_/C _13736_/X vssd1 vssd1 vccd1 vccd1 _13899_/Y sky130_fd_sc_hd__a21oi_1
X_16687_ _16687_/A _07784_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16630__35 vssd1 vssd1 vccd1 vccd1 _16630__35/HI _16696_/A sky130_fd_sc_hd__conb_1
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15638_ _15791_/CLK _15638_/D vssd1 vssd1 vccd1 vccd1 _15638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _16551_/CLK _15569_/D vssd1 vssd1 vccd1 vccd1 _15569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _08110_/A vssd1 vssd1 vccd1 vccd1 _08766_/C sky130_fd_sc_hd__clkbuf_2
X_09090_ _09756_/A vssd1 vssd1 vccd1 vccd1 _09090_/X sky130_fd_sc_hd__clkbuf_2
X_08041_ _16433_/Q vssd1 vssd1 vccd1 vccd1 _14559_/A sky130_fd_sc_hd__clkinv_2
XFILLER_128_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09992_ _15737_/Q _09992_/B _09998_/C vssd1 vssd1 vccd1 vccd1 _09994_/C sky130_fd_sc_hd__nand3_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ _15523_/Q _08943_/B _08948_/C vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__and3_1
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08874_ _08916_/A _08880_/C vssd1 vssd1 vccd1 vccd1 _08874_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07825_ _07837_/A vssd1 vssd1 vccd1 vccd1 _07830_/A sky130_fd_sc_hd__buf_12
X_07756_ input1/X vssd1 vssd1 vccd1 vccd1 _07849_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09426_ _09423_/A _09423_/B _09422_/Y _09425_/Y vssd1 vssd1 vccd1 vccd1 _15619_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09357_ _09360_/C vssd1 vssd1 vccd1 vccd1 _09371_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08308_ _15448_/Q _08415_/A vssd1 vssd1 vccd1 vccd1 _08309_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09288_ _09286_/X _09288_/B vssd1 vssd1 vccd1 vccd1 _09288_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08239_ _14559_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08239_/X sky130_fd_sc_hd__or2_1
XFILLER_125_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11250_ _11250_/A vssd1 vssd1 vccd1 vccd1 _15944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10201_ _10250_/A _10201_/B _10201_/C vssd1 vssd1 vccd1 vccd1 _10202_/A sky130_fd_sc_hd__and3_1
XFILLER_106_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11181_ _12029_/A vssd1 vssd1 vccd1 vccd1 _11181_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10132_ _15764_/Q _10133_/C _09813_/X vssd1 vssd1 vccd1 vccd1 _10132_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10063_ _10061_/A _10061_/B _10062_/X vssd1 vssd1 vccd1 vccd1 _15747_/D sky130_fd_sc_hd__a21oi_1
XFILLER_88_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14940_ _16476_/Q _14995_/B _14940_/C vssd1 vssd1 vccd1 vccd1 _14949_/A sky130_fd_sc_hd__and3_1
XFILLER_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14871_ _14871_/A vssd1 vssd1 vccd1 vccd1 _16464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16610_ input11/X _16610_/D vssd1 vssd1 vccd1 vccd1 _16610_/Q sky130_fd_sc_hd__dfxtp_1
X_13822_ _16309_/Q _13929_/B _13822_/C vssd1 vssd1 vccd1 vccd1 _13831_/B sky130_fd_sc_hd__and3_1
XFILLER_29_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ _16595_/CLK _16541_/D vssd1 vssd1 vccd1 vccd1 _16710_/A sky130_fd_sc_hd__dfxtp_1
X_13753_ _16298_/Q _13753_/B _13759_/C vssd1 vssd1 vccd1 vccd1 _13753_/Y sky130_fd_sc_hd__nand3_1
XFILLER_141_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10965_ _10959_/C _10960_/C _10962_/Y _10963_/X vssd1 vssd1 vccd1 vccd1 _10966_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ _12704_/A vssd1 vssd1 vccd1 vccd1 _12718_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16472_ input11/X _16472_/D vssd1 vssd1 vccd1 vccd1 _16472_/Q sky130_fd_sc_hd__dfxtp_1
X_13684_ _16289_/Q _13856_/B _13684_/C vssd1 vssd1 vccd1 vccd1 _13684_/Y sky130_fd_sc_hd__nand3_1
X_10896_ _10954_/A _10896_/B _10902_/A vssd1 vssd1 vccd1 vccd1 _15894_/D sky130_fd_sc_hd__nor3_1
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15423_ _16237_/Q _16236_/Q _16235_/Q _15422_/X vssd1 vssd1 vccd1 vccd1 _16600_/D
+ sky130_fd_sc_hd__o31a_1
X_12635_ _12635_/A _12643_/B vssd1 vssd1 vccd1 vccd1 _12637_/A sky130_fd_sc_hd__or2_1
XFILLER_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15354_ _09076_/A _15347_/B _15350_/B _15353_/Y vssd1 vssd1 vccd1 vccd1 _16548_/D
+ sky130_fd_sc_hd__o31a_1
X_12566_ _12566_/A vssd1 vssd1 vccd1 vccd1 _16130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11517_ _12650_/A vssd1 vssd1 vccd1 vccd1 _11517_/X sky130_fd_sc_hd__clkbuf_2
X_14305_ _14303_/Y _14299_/C _14301_/Y _14302_/X vssd1 vssd1 vccd1 vccd1 _14306_/C
+ sky130_fd_sc_hd__a211o_1
X_15285_ _16706_/A _15306_/A vssd1 vssd1 vccd1 vccd1 _15286_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _12495_/Y _12490_/C _12492_/Y _12493_/X vssd1 vssd1 vccd1 vccd1 _12498_/C
+ sky130_fd_sc_hd__a211o_1
X_14236_ _14799_/A vssd1 vssd1 vccd1 vccd1 _14458_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_11448_ _11617_/A _11452_/C vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__or2_1
XFILLER_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ _14187_/C vssd1 vssd1 vccd1 vccd1 _14201_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11379_ _11379_/A _11379_/B _11383_/B vssd1 vssd1 vccd1 vccd1 _15963_/D sky130_fd_sc_hd__nor3_1
XFILLER_140_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13682_/A vssd1 vssd1 vccd1 vccd1 _13342_/B sky130_fd_sc_hd__clkbuf_2
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14096_/Y _14090_/C _14093_/Y _14103_/A vssd1 vssd1 vccd1 vccd1 _14103_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13049_ _13049_/A _13049_/B _13049_/C vssd1 vssd1 vccd1 vccd1 _13050_/C sky130_fd_sc_hd__nand3_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08590_ _15459_/Q _08807_/B _08590_/C vssd1 vssd1 vccd1 vccd1 _08592_/C sky130_fd_sc_hd__nand3_1
XFILLER_54_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16739_ _16739_/A _07846_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09211_ _09220_/C vssd1 vssd1 vccd1 vccd1 _09231_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09142_ _09142_/A _09142_/B _09142_/C vssd1 vssd1 vccd1 vccd1 _09143_/A sky130_fd_sc_hd__and3_1
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09073_ _09073_/A _09073_/B vssd1 vssd1 vccd1 vccd1 _09074_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08024_ _16562_/Q vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__inv_2
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09975_ _09307_/X _09973_/B _09894_/X vssd1 vssd1 vccd1 vccd1 _09975_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08926_ _08926_/A _08926_/B vssd1 vssd1 vccd1 vccd1 _15514_/D sky130_fd_sc_hd__nor2_1
XFILLER_130_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08857_ _10782_/B vssd1 vssd1 vccd1 vccd1 _10492_/A sky130_fd_sc_hd__buf_4
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07808_ _07811_/A vssd1 vssd1 vccd1 vccd1 _07808_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08788_ _08831_/A _08791_/C vssd1 vssd1 vccd1 vccd1 _08790_/A sky130_fd_sc_hd__and2_1
XFILLER_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10750_ _15873_/Q _10750_/B _10755_/C vssd1 vssd1 vccd1 vccd1 _10750_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09409_ _09629_/A vssd1 vssd1 vccd1 vccd1 _09585_/B sky130_fd_sc_hd__buf_2
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ _10681_/A _10681_/B _10681_/C vssd1 vssd1 vccd1 vccd1 _10682_/C sky130_fd_sc_hd__nand3_1
XFILLER_41_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _12420_/A vssd1 vssd1 vccd1 vccd1 _16109_/D sky130_fd_sc_hd__clkbuf_1
X_12351_ _16101_/Q _12352_/C _12292_/X vssd1 vssd1 vccd1 vccd1 _12353_/A sky130_fd_sc_hd__a21oi_1
XFILLER_138_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ _11300_/Y _11301_/X _11297_/C _11298_/C vssd1 vssd1 vccd1 vccd1 _11304_/B
+ sky130_fd_sc_hd__o211ai_1
X_15070_ _15083_/C vssd1 vssd1 vccd1 vccd1 _15090_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12282_ _12280_/Y _12274_/C _12276_/Y _12279_/X vssd1 vssd1 vccd1 vccd1 _12283_/C
+ sky130_fd_sc_hd__a211o_1
X_14021_ _14021_/A vssd1 vssd1 vccd1 vccd1 _16336_/D sky130_fd_sc_hd__clkbuf_1
X_11233_ _11233_/A vssd1 vssd1 vccd1 vccd1 _11233_/X sky130_fd_sc_hd__buf_4
XFILLER_107_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11164_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11169_/C sky130_fd_sc_hd__nor2_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10115_ _09851_/X _10107_/B _10110_/B _10114_/Y vssd1 vssd1 vccd1 vccd1 _15757_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15972_ _16005_/CLK _15972_/D vssd1 vssd1 vccd1 vccd1 _15972_/Q sky130_fd_sc_hd__dfxtp_1
X_11095_ _11090_/Y _11101_/A _11094_/Y _11088_/C vssd1 vssd1 vccd1 vccd1 _11097_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10046_ _10043_/Y _10044_/X _10045_/Y _10041_/C vssd1 vssd1 vccd1 vccd1 _10048_/B
+ sky130_fd_sc_hd__o211ai_1
X_14923_ _16474_/Q _14925_/C _14694_/X vssd1 vssd1 vccd1 vccd1 _14923_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14854_ _14855_/B _14855_/C _14855_/A vssd1 vssd1 vccd1 vccd1 _14856_/B sky130_fd_sc_hd__a21o_1
XFILLER_17_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13805_ _16307_/Q _13815_/C _13750_/X vssd1 vssd1 vccd1 vccd1 _13805_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11997_ _11995_/Y _11990_/C _11992_/Y _11994_/X vssd1 vssd1 vccd1 vccd1 _11998_/C
+ sky130_fd_sc_hd__a211o_1
X_14785_ _14785_/A vssd1 vssd1 vccd1 vccd1 _14800_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16524_ _16595_/CLK _16524_/D vssd1 vssd1 vccd1 vccd1 _16524_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10948_ _10963_/C vssd1 vssd1 vccd1 vccd1 _10970_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13736_ _14015_/A vssd1 vssd1 vccd1 vccd1 _13736_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16455_ input11/X _16455_/D vssd1 vssd1 vccd1 vccd1 _16455_/Q sky130_fd_sc_hd__dfxtp_1
X_13667_ _16288_/Q _13676_/C _13443_/X vssd1 vssd1 vccd1 vccd1 _13670_/B sky130_fd_sc_hd__a21o_1
X_10879_ _10879_/A _10886_/B vssd1 vssd1 vccd1 vccd1 _10881_/A sky130_fd_sc_hd__or2_1
X_15406_ _16133_/Q _16132_/Q _16131_/Q _15403_/X vssd1 vssd1 vccd1 vccd1 _16587_/D
+ sky130_fd_sc_hd__o31a_1
X_12618_ _12618_/A vssd1 vssd1 vccd1 vccd1 _16137_/D sky130_fd_sc_hd__clkbuf_1
X_16386_ _16389_/CLK _16386_/D vssd1 vssd1 vccd1 vccd1 _16386_/Q sky130_fd_sc_hd__dfxtp_1
X_13598_ _13598_/A vssd1 vssd1 vccd1 vccd1 _13635_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12549_ _12549_/A vssd1 vssd1 vccd1 vccd1 _16128_/D sky130_fd_sc_hd__clkbuf_1
X_15337_ _15337_/A _15337_/B _15337_/C vssd1 vssd1 vccd1 vccd1 _15338_/C sky130_fd_sc_hd__nand3_1
XFILLER_129_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _07824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15268_ _15268_/A _15274_/B vssd1 vssd1 vccd1 vccd1 _15270_/A sky130_fd_sc_hd__or2_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14219_ _14219_/A vssd1 vssd1 vccd1 vccd1 _16365_/D sky130_fd_sc_hd__clkbuf_1
X_15199_ _15199_/A vssd1 vssd1 vccd1 vccd1 _16518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _15691_/Q _09781_/C _09714_/X vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__a21oi_1
XFILLER_140_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08711_ _15350_/A vssd1 vssd1 vccd1 vccd1 _08711_/X sky130_fd_sc_hd__clkbuf_2
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09691_ _09688_/A _09687_/Y _09688_/B vssd1 vssd1 vccd1 vccd1 _09691_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08642_ _08831_/A _08651_/C vssd1 vssd1 vccd1 vccd1 _08646_/A sky130_fd_sc_hd__and2_1
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _09801_/A vssd1 vssd1 vccd1 vccd1 _12932_/A sky130_fd_sc_hd__buf_6
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ _09125_/A vssd1 vssd1 vccd1 vccd1 _09125_/X sky130_fd_sc_hd__clkbuf_2
X_09056_ _09056_/A vssd1 vssd1 vccd1 vccd1 _09220_/B sky130_fd_sc_hd__buf_2
X_08007_ _16584_/Q vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__inv_2
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09958_ _10055_/A _09958_/B _09961_/B vssd1 vssd1 vccd1 vccd1 _15726_/D sky130_fd_sc_hd__nor3_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16666__71 vssd1 vssd1 vccd1 vccd1 _16666__71/HI _16742_/A sky130_fd_sc_hd__conb_1
XFILLER_58_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08909_ _08909_/A _08909_/B vssd1 vssd1 vccd1 vccd1 _08911_/B sky130_fd_sc_hd__nor2_1
X_09889_ _09883_/Y _09884_/X _09886_/B vssd1 vssd1 vccd1 vccd1 _09890_/B sky130_fd_sc_hd__o21a_1
XFILLER_58_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ _11920_/A vssd1 vssd1 vccd1 vccd1 _16039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11851_ _11852_/B _11852_/C _11850_/X vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__o21ai_1
XFILLER_73_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10802_ _10802_/A vssd1 vssd1 vccd1 vccd1 _15881_/D sky130_fd_sc_hd__clkbuf_1
X_14570_ _14571_/B _14571_/C _14571_/A vssd1 vssd1 vccd1 vccd1 _14572_/B sky130_fd_sc_hd__a21o_1
X_11782_ _11780_/Y _11776_/C _11778_/Y _11787_/A vssd1 vssd1 vccd1 vccd1 _11787_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_26_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _10733_/A vssd1 vssd1 vccd1 vccd1 _15869_/D sky130_fd_sc_hd__clkbuf_1
X_13521_ _13521_/A vssd1 vssd1 vccd1 vccd1 _14647_/A sky130_fd_sc_hd__clkbuf_8
X_16240_ _16261_/CLK _16240_/D vssd1 vssd1 vccd1 vccd1 _16240_/Q sky130_fd_sc_hd__dfxtp_1
X_13452_ _16257_/Q _13617_/B _13452_/C vssd1 vssd1 vccd1 vccd1 _13452_/X sky130_fd_sc_hd__and3_1
XFILLER_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10664_ _10659_/B _10662_/B _08705_/B vssd1 vssd1 vccd1 vccd1 _10665_/B sky130_fd_sc_hd__o21a_1
X_12403_ _12686_/A vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__clkbuf_2
X_13383_ _16247_/Q _13383_/B _13393_/C vssd1 vssd1 vccd1 vccd1 _13388_/A sky130_fd_sc_hd__and3_1
X_16171_ _16237_/CLK _16171_/D vssd1 vssd1 vccd1 vccd1 _16171_/Q sky130_fd_sc_hd__dfxtp_1
X_10595_ _10588_/C _10589_/C _10592_/Y _10593_/X vssd1 vssd1 vccd1 vccd1 _10596_/C
+ sky130_fd_sc_hd__a211o_1
X_15122_ _15135_/C vssd1 vssd1 vccd1 vccd1 _15142_/C sky130_fd_sc_hd__clkbuf_1
X_12334_ _12332_/Y _12328_/C _12330_/Y _12331_/X vssd1 vssd1 vccd1 vccd1 _12335_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15053_ _15053_/A _15053_/B _15057_/B vssd1 vssd1 vccd1 vccd1 _16493_/D sky130_fd_sc_hd__nor3_1
X_12265_ _12257_/C _12258_/C _12260_/Y _12263_/X vssd1 vssd1 vccd1 vccd1 _12266_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14004_ _16335_/Q _14044_/C _13781_/X vssd1 vssd1 vccd1 vccd1 _14007_/B sky130_fd_sc_hd__a21oi_1
X_11216_ _15941_/Q _11217_/C _11158_/X vssd1 vssd1 vccd1 vccd1 _11218_/A sky130_fd_sc_hd__a21oi_1
X_12196_ _12230_/A _12196_/B _12200_/A vssd1 vssd1 vccd1 vccd1 _16078_/D sky130_fd_sc_hd__nor3_1
XFILLER_96_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11147_ _11145_/Y _11140_/C _11142_/Y _11144_/X vssd1 vssd1 vccd1 vccd1 _11148_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15955_ _15365_/A _15955_/D vssd1 vssd1 vccd1 vccd1 _15955_/Q sky130_fd_sc_hd__dfxtp_1
X_11078_ _15921_/Q _11309_/B _11078_/C vssd1 vssd1 vccd1 vccd1 _11078_/Y sky130_fd_sc_hd__nand3_1
XFILLER_76_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10029_ _15744_/Q _10178_/B _10029_/C vssd1 vssd1 vccd1 vccd1 _10034_/A sky130_fd_sc_hd__and3_1
X_14906_ _14906_/A vssd1 vssd1 vccd1 vccd1 _14906_/X sky130_fd_sc_hd__clkbuf_2
X_15886_ _16553_/Q _15886_/D vssd1 vssd1 vccd1 vccd1 _15886_/Q sky130_fd_sc_hd__dfxtp_2
X_14837_ _15007_/A vssd1 vssd1 vccd1 vccd1 _14878_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14768_ _14768_/A _14768_/B _14772_/B vssd1 vssd1 vccd1 vccd1 _16448_/D sky130_fd_sc_hd__nor3_1
X_16507_ _16607_/CLK _16507_/D vssd1 vssd1 vccd1 vccd1 _16507_/Q sky130_fd_sc_hd__dfxtp_1
X_13719_ _13719_/A vssd1 vssd1 vccd1 vccd1 _16293_/D sky130_fd_sc_hd__clkbuf_1
X_14699_ _14697_/Y _14692_/C _14695_/Y _14696_/X vssd1 vssd1 vccd1 vccd1 _14700_/C
+ sky130_fd_sc_hd__a211o_1
X_16438_ _16595_/CLK _16438_/D vssd1 vssd1 vccd1 vccd1 _16438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16369_ _16389_/CLK _16369_/D vssd1 vssd1 vccd1 vccd1 _16369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09812_ _09812_/A vssd1 vssd1 vccd1 vccd1 _09951_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ _09737_/Y _09741_/X _09742_/Y vssd1 vssd1 vccd1 vccd1 _15683_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09674_ _09674_/A _09674_/B _09674_/C vssd1 vssd1 vccd1 vccd1 _09675_/C sky130_fd_sc_hd__nand3_1
XFILLER_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ input4/X vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__buf_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08556_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08556_/X sky130_fd_sc_hd__and2_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08487_ _08487_/A _08487_/B vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ _09148_/A _09108_/B _09112_/B vssd1 vssd1 vccd1 vccd1 _15555_/D sky130_fd_sc_hd__nor3_1
XFILLER_109_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10380_ _10429_/A _10380_/B _10384_/A vssd1 vssd1 vccd1 vccd1 _15805_/D sky130_fd_sc_hd__nor3_1
XFILLER_136_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09039_ _09126_/A vssd1 vssd1 vccd1 vccd1 _09039_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ _12901_/A vssd1 vssd1 vccd1 vccd1 _12050_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11001_ _11169_/A _11001_/B _11001_/C vssd1 vssd1 vccd1 vccd1 _11002_/C sky130_fd_sc_hd__or3_1
XFILLER_132_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15740_ _15812_/CLK _15740_/D vssd1 vssd1 vccd1 vccd1 _15740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12952_ _16185_/Q _13009_/B _12952_/C vssd1 vssd1 vccd1 vccd1 _12952_/Y sky130_fd_sc_hd__nand3_1
XFILLER_133_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11903_ _11903_/A vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _15791_/CLK _15671_/D vssd1 vssd1 vccd1 vccd1 _15671_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12883_ _12883_/A _12883_/B _12883_/C vssd1 vssd1 vccd1 vccd1 _12884_/C sky130_fd_sc_hd__nand3_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _16426_/Q _14662_/C _14621_/X vssd1 vssd1 vccd1 vccd1 _14624_/B sky130_fd_sc_hd__a21oi_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _11963_/A vssd1 vssd1 vccd1 vccd1 _11948_/A sky130_fd_sc_hd__buf_2
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11765_ _11762_/Y _11763_/X _11764_/Y _11760_/C vssd1 vssd1 vccd1 vccd1 _11767_/B
+ sky130_fd_sc_hd__o211ai_1
X_14553_ _14722_/A vssd1 vssd1 vccd1 vccd1 _14594_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _13526_/A _13504_/B _13504_/C vssd1 vssd1 vccd1 vccd1 _13505_/A sky130_fd_sc_hd__and3_1
X_10716_ _10716_/A vssd1 vssd1 vccd1 vccd1 _10716_/X sky130_fd_sc_hd__buf_2
XFILLER_147_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11696_ _16009_/Q _11706_/C _11471_/X vssd1 vssd1 vccd1 vccd1 _11696_/Y sky130_fd_sc_hd__a21oi_1
X_14484_ _14484_/A _14484_/B _14488_/B vssd1 vssd1 vccd1 vccd1 _16403_/D sky130_fd_sc_hd__nor3_1
X_16223_ _16261_/CLK _16223_/D vssd1 vssd1 vccd1 vccd1 _16223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ _10644_/Y _10645_/X _10646_/Y _10642_/C vssd1 vssd1 vccd1 vccd1 _10649_/B
+ sky130_fd_sc_hd__o211ai_1
X_13435_ _13435_/A vssd1 vssd1 vccd1 vccd1 _13452_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16154_ _16555_/Q _16154_/D vssd1 vssd1 vccd1 vccd1 _16154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13366_ _13366_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__nor2_1
X_10578_ _10578_/A vssd1 vssd1 vccd1 vccd1 _10676_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105_ _15102_/Y _15111_/A _15104_/Y _15100_/C vssd1 vssd1 vccd1 vccd1 _15107_/B
+ sky130_fd_sc_hd__o211a_1
X_12317_ _16096_/Q _12325_/C _12316_/X vssd1 vssd1 vccd1 vccd1 _12320_/B sky130_fd_sc_hd__a21o_1
X_16085_ _16554_/Q _16085_/D vssd1 vssd1 vccd1 vccd1 _16085_/Q sky130_fd_sc_hd__dfxtp_1
X_13297_ _16235_/Q _13305_/C _13184_/X vssd1 vssd1 vccd1 vccd1 _13297_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12248_ _12263_/C vssd1 vssd1 vccd1 vccd1 _12271_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15036_ _15032_/Y _15033_/X _15035_/Y _15030_/C vssd1 vssd1 vccd1 vccd1 _15038_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_69_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12179_ _16077_/Q _12232_/B _12179_/C vssd1 vssd1 vccd1 vccd1 _12187_/B sky130_fd_sc_hd__and3_1
XFILLER_122_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15938_ _15365_/A _15938_/D vssd1 vssd1 vccd1 vccd1 _15938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15869_ _16570_/CLK _15869_/D vssd1 vssd1 vccd1 vccd1 _15869_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08410_ _08410_/A _08410_/B vssd1 vssd1 vccd1 vccd1 _08431_/A sky130_fd_sc_hd__xnor2_1
X_09390_ _09436_/A _09390_/B vssd1 vssd1 vccd1 vccd1 _09390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08341_ _08139_/A _08139_/B _08340_/X vssd1 vssd1 vccd1 vccd1 _08435_/B sky130_fd_sc_hd__a21oi_4
X_08272_ _08273_/A _08273_/B vssd1 vssd1 vccd1 vccd1 _08274_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07987_ _08186_/B _07987_/B vssd1 vssd1 vccd1 vccd1 _08004_/A sky130_fd_sc_hd__nand2_2
X_16636__41 vssd1 vssd1 vccd1 vccd1 _16636__41/HI _16712_/A sky130_fd_sc_hd__conb_1
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09726_ _15684_/Q _09727_/C _09590_/X vssd1 vssd1 vccd1 vccd1 _09726_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09657_ _09524_/X _09655_/B _09656_/Y vssd1 vssd1 vccd1 vccd1 _15666_/D sky130_fd_sc_hd__o21a_1
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08608_ _15460_/Q _10743_/B _08619_/C vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__and3_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09588_ _09588_/A _09588_/B _09588_/C vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__and3_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08540_/B _08540_/C _08540_/A vssd1 vssd1 vccd1 vccd1 _08541_/A sky130_fd_sc_hd__a21oi_1
XFILLER_70_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11550_ _15988_/Q _11560_/C _11434_/X vssd1 vssd1 vccd1 vccd1 _11550_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ _10501_/A vssd1 vssd1 vccd1 vccd1 _10691_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ _11478_/Y _11479_/X _11480_/Y _11476_/C vssd1 vssd1 vccd1 vccd1 _11483_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13220_ _16224_/Q _13228_/C _13162_/X vssd1 vssd1 vccd1 vccd1 _13224_/B sky130_fd_sc_hd__a21o_1
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10432_ _10486_/A vssd1 vssd1 vccd1 vccd1 _10432_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13151_ _13151_/A _13151_/B _13151_/C vssd1 vssd1 vccd1 vccd1 _13152_/C sky130_fd_sc_hd__or3_1
X_10363_ _10363_/A _10363_/B vssd1 vssd1 vccd1 vccd1 _10365_/A sky130_fd_sc_hd__or2_1
X_12102_ _12100_/Y _12096_/C _12098_/Y _12099_/X vssd1 vssd1 vccd1 vccd1 _12103_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13082_ _16205_/Q _13082_/B _13082_/C vssd1 vssd1 vccd1 vccd1 _13093_/B sky130_fd_sc_hd__and3_1
X_10294_ _15791_/Q _10294_/B _10294_/C vssd1 vssd1 vccd1 vccd1 _10294_/X sky130_fd_sc_hd__and3_1
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12033_ _12033_/A _12033_/B _12033_/C vssd1 vssd1 vccd1 vccd1 _12034_/C sky130_fd_sc_hd__nand3_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13984_ _13982_/Y _13977_/C _13980_/Y _13991_/A vssd1 vssd1 vccd1 vccd1 _13991_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_92_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15723_ _15812_/CLK _15723_/D vssd1 vssd1 vccd1 vccd1 _15723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12935_ _16183_/Q _13102_/B _12945_/C vssd1 vssd1 vccd1 vccd1 _12941_/A sky130_fd_sc_hd__and3_1
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15654_ _15791_/CLK _15654_/D vssd1 vssd1 vccd1 vccd1 _15654_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _13034_/A vssd1 vssd1 vccd1 vccd1 _12907_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _14605_/A _14605_/B vssd1 vssd1 vccd1 vccd1 _14606_/B sky130_fd_sc_hd__nor2_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _11832_/A _11817_/B _11817_/C vssd1 vssd1 vccd1 vccd1 _11818_/A sky130_fd_sc_hd__and3_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _16551_/CLK _15585_/D vssd1 vssd1 vccd1 vccd1 _15585_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _16165_/Q _12798_/C _12575_/X vssd1 vssd1 vccd1 vccd1 _12799_/A sky130_fd_sc_hd__a21oi_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _14536_/A vssd1 vssd1 vccd1 vccd1 _16411_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _12029_/A vssd1 vssd1 vccd1 vccd1 _11748_/X sky130_fd_sc_hd__clkbuf_2
X_14467_ _14463_/Y _14464_/X _14466_/Y _14461_/C vssd1 vssd1 vccd1 vccd1 _14469_/B
+ sky130_fd_sc_hd__o211ai_1
X_11679_ _11737_/A _11679_/B _11679_/C vssd1 vssd1 vccd1 vccd1 _11680_/C sky130_fd_sc_hd__or3_1
X_16206_ _16237_/CLK _16206_/D vssd1 vssd1 vccd1 vccd1 _16206_/Q sky130_fd_sc_hd__dfxtp_2
X_13418_ _13415_/Y _13426_/A _13417_/Y _13412_/C vssd1 vssd1 vccd1 vccd1 _13420_/B
+ sky130_fd_sc_hd__o211a_1
X_14398_ _14484_/A _14398_/B _14402_/A vssd1 vssd1 vccd1 vccd1 _16390_/D sky130_fd_sc_hd__nor3_1
XFILLER_143_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _16555_/Q _16137_/D vssd1 vssd1 vccd1 vccd1 _16137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13349_ _16243_/Q _13358_/C _13184_/X vssd1 vssd1 vccd1 vccd1 _13349_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16068_ _16554_/Q _16068_/D vssd1 vssd1 vccd1 vccd1 _16068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15019_ _15053_/A _15019_/B _15023_/A vssd1 vssd1 vccd1 vccd1 _16488_/D sky130_fd_sc_hd__nor3_1
X_07910_ _07910_/A _07910_/B vssd1 vssd1 vccd1 vccd1 _07911_/B sky130_fd_sc_hd__nand2_2
X_08890_ _08896_/C vssd1 vssd1 vccd1 vccd1 _08907_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07841_ _07842_/A vssd1 vssd1 vccd1 vccd1 _07841_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07772_ _07774_/A vssd1 vssd1 vccd1 vccd1 _07772_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ _15640_/Q _09519_/C _09463_/X vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__a21oi_1
XFILLER_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09442_ _09396_/X _10526_/A _09436_/B _08554_/A vssd1 vssd1 vccd1 vccd1 _09443_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _09366_/C _09367_/C _09370_/Y _09377_/A vssd1 vssd1 vccd1 vccd1 _09377_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_40_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08324_ _08195_/A _08195_/B _08323_/X vssd1 vssd1 vccd1 vccd1 _08344_/A sky130_fd_sc_hd__a21bo_1
X_08255_ _08978_/C _08083_/B _08082_/B vssd1 vssd1 vccd1 vccd1 _08259_/A sky130_fd_sc_hd__o21a_1
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08186_ _08186_/A _08186_/B _08186_/C vssd1 vssd1 vccd1 vccd1 _08187_/B sky130_fd_sc_hd__nand3_1
XFILLER_146_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _09709_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _15677_/D sky130_fd_sc_hd__nor2_1
XFILLER_74_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10981_ _10981_/A _10981_/B _10981_/C vssd1 vssd1 vccd1 vccd1 _10982_/A sky130_fd_sc_hd__and3_1
X_12720_ _12714_/C _12715_/C _12717_/Y _12718_/X vssd1 vssd1 vccd1 vccd1 _12721_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12651_ _16143_/Q _12692_/C _12650_/X vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__a21oi_1
XFILLER_71_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11602_ _11599_/Y _11600_/X _11601_/Y _11597_/C vssd1 vssd1 vccd1 vccd1 _11604_/B
+ sky130_fd_sc_hd__o211ai_1
X_15370_ _15901_/Q _15900_/Q _15899_/Q _15363_/X vssd1 vssd1 vccd1 vccd1 _16558_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12582_ _12749_/A _12586_/C vssd1 vssd1 vccd1 vccd1 _12582_/X sky130_fd_sc_hd__or2_1
XFILLER_90_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14321_ _14342_/A _14321_/B _14325_/B vssd1 vssd1 vccd1 vccd1 _16379_/D sky130_fd_sc_hd__nor3_1
X_11533_ _11533_/A vssd1 vssd1 vccd1 vccd1 _15984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ _15976_/Q _11473_/C _11463_/X vssd1 vssd1 vccd1 vccd1 _11467_/B sky130_fd_sc_hd__a21o_1
X_14252_ _16371_/Q _14472_/B _14260_/C vssd1 vssd1 vccd1 vccd1 _14252_/X sky130_fd_sc_hd__and3_1
XFILLER_109_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ _10409_/B _10412_/B _10414_/X vssd1 vssd1 vccd1 vccd1 _10416_/B sky130_fd_sc_hd__o21a_1
X_13203_ _13315_/A _13209_/C vssd1 vssd1 vccd1 vccd1 _13203_/X sky130_fd_sc_hd__or2_1
X_11395_ _14220_/A vssd1 vssd1 vccd1 vccd1 _11963_/A sky130_fd_sc_hd__buf_2
X_14183_ _14183_/A vssd1 vssd1 vccd1 vccd1 _16360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10346_ _10346_/A vssd1 vssd1 vccd1 vccd1 _15798_/D sky130_fd_sc_hd__clkbuf_1
X_13134_ _16212_/Q _13143_/C _13133_/X vssd1 vssd1 vccd1 vccd1 _13134_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13072_/A _13065_/B _13065_/C vssd1 vssd1 vccd1 vccd1 _13066_/A sky130_fd_sc_hd__and3_1
XFILLER_124_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10277_ _10168_/X _10274_/B _10224_/X vssd1 vssd1 vccd1 vccd1 _10277_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12016_ _12185_/A vssd1 vssd1 vccd1 vccd1 _12056_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16755_ _16755_/A _07773_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
XFILLER_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13967_ _13963_/Y _13965_/X _13966_/Y _13961_/C vssd1 vssd1 vccd1 vccd1 _13969_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15706_ _15812_/CLK _15706_/D vssd1 vssd1 vccd1 vccd1 _15706_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12918_ _12918_/A _12918_/B vssd1 vssd1 vccd1 vccd1 _12919_/B sky130_fd_sc_hd__nor2_1
X_16686_ _16686_/A _07783_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13898_ _13898_/A vssd1 vssd1 vccd1 vccd1 _16319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15637_ _15791_/CLK _15637_/D vssd1 vssd1 vccd1 vccd1 _15637_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _12849_/A vssd1 vssd1 vccd1 vccd1 _13979_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15568_ _16551_/CLK _15568_/D vssd1 vssd1 vccd1 vccd1 _15568_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14519_ _14535_/A _14519_/B _14519_/C vssd1 vssd1 vccd1 vccd1 _14520_/A sky130_fd_sc_hd__and3_1
X_15499_ _16570_/CLK _15499_/D vssd1 vssd1 vccd1 vccd1 _15499_/Q sky130_fd_sc_hd__dfxtp_2
X_08040_ _16586_/Q vssd1 vssd1 vccd1 vccd1 _12473_/A sky130_fd_sc_hd__clkinv_4
XFILLER_116_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09991_ _15737_/Q _09998_/C _08589_/A vssd1 vssd1 vccd1 vccd1 _09994_/B sky130_fd_sc_hd__a21o_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ _15523_/Q _08948_/C _08859_/X vssd1 vssd1 vccd1 vccd1 _08942_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08873_ _08867_/B _08870_/B _08698_/X vssd1 vssd1 vccd1 vccd1 _08880_/C sky130_fd_sc_hd__o21a_1
XFILLER_97_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07824_ _07824_/A vssd1 vssd1 vccd1 vccd1 _07824_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09425_ _09423_/X _09422_/Y _09424_/X vssd1 vssd1 vccd1 vccd1 _09425_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _15624_/Q vssd1 vssd1 vccd1 vccd1 _09360_/C sky130_fd_sc_hd__inv_2
X_08307_ _16703_/A vssd1 vssd1 vccd1 vccd1 _08415_/A sky130_fd_sc_hd__inv_2
XFILLER_138_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09287_ _15596_/Q _09286_/C _09117_/A vssd1 vssd1 vccd1 vccd1 _09288_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08238_ _08383_/A _08238_/B vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__nand2_2
XFILLER_107_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08169_ _08169_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08171_/B sky130_fd_sc_hd__xnor2_1
XFILLER_109_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10200_ _10198_/Y _10193_/C _10195_/Y _10197_/X vssd1 vssd1 vccd1 vccd1 _10201_/C
+ sky130_fd_sc_hd__a211o_1
X_11180_ _11236_/A _11180_/B _11185_/A vssd1 vssd1 vccd1 vccd1 _15934_/D sky130_fd_sc_hd__nor3_1
XFILLER_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10131_ _10131_/A vssd1 vssd1 vccd1 vccd1 _15761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _10271_/A _10062_/B vssd1 vssd1 vccd1 vccd1 _10062_/X sky130_fd_sc_hd__or2_1
XFILLER_125_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14870_ _14878_/A _14870_/B _14870_/C vssd1 vssd1 vccd1 vccd1 _14871_/A sky130_fd_sc_hd__and3_1
X_13821_ _16309_/Q _13822_/C _13705_/X vssd1 vssd1 vccd1 vccd1 _13823_/A sky130_fd_sc_hd__a21oi_1
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16540_ _16595_/CLK _16540_/D vssd1 vssd1 vccd1 vccd1 _16709_/A sky130_fd_sc_hd__dfxtp_1
X_13752_ _16299_/Q _13914_/B _13759_/C vssd1 vssd1 vccd1 vccd1 _13752_/X sky130_fd_sc_hd__and3_1
X_10964_ _10962_/Y _10963_/X _10959_/C _10960_/C vssd1 vssd1 vccd1 vccd1 _10966_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12703_ _12703_/A vssd1 vssd1 vccd1 vccd1 _16149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16471_ _16607_/CLK _16471_/D vssd1 vssd1 vccd1 vccd1 _16471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13683_ _16290_/Q _13906_/B _13684_/C vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__and3_1
XFILLER_71_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10895_ _15895_/Q _11118_/B _10907_/C vssd1 vssd1 vccd1 vccd1 _10902_/A sky130_fd_sc_hd__and3_1
X_15422_ _15440_/A vssd1 vssd1 vccd1 vccd1 _15422_/X sky130_fd_sc_hd__clkbuf_2
X_12634_ _16141_/Q _12798_/B _12634_/C vssd1 vssd1 vccd1 vccd1 _12643_/B sky130_fd_sc_hd__and3_1
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15353_ _15353_/A _15358_/C vssd1 vssd1 vccd1 vccd1 _15353_/Y sky130_fd_sc_hd__nor2_1
X_12565_ _12565_/A _12565_/B _12565_/C vssd1 vssd1 vccd1 vccd1 _12566_/A sky130_fd_sc_hd__and3_1
XFILLER_12_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ _14301_/Y _14302_/X _14303_/Y _14299_/C vssd1 vssd1 vccd1 vccd1 _14306_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_129_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ _12932_/A vssd1 vssd1 vccd1 vccd1 _12650_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15284_ _16702_/A vssd1 vssd1 vccd1 vccd1 _15306_/A sky130_fd_sc_hd__inv_2
X_12496_ _12492_/Y _12493_/X _12495_/Y _12490_/C vssd1 vssd1 vccd1 vccd1 _12498_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_116_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14235_ _16369_/Q _14245_/C _14015_/X vssd1 vssd1 vccd1 vccd1 _14235_/Y sky130_fd_sc_hd__a21oi_1
X_11447_ _11447_/A _11447_/B vssd1 vssd1 vccd1 vccd1 _11452_/C sky130_fd_sc_hd__nor2_1
XFILLER_137_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11378_ _11376_/Y _11371_/C _11373_/Y _11383_/A vssd1 vssd1 vccd1 vccd1 _11383_/B
+ sky130_fd_sc_hd__a211oi_1
X_14166_ _14179_/C vssd1 vssd1 vccd1 vccd1 _14187_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _10342_/C vssd1 vssd1 vccd1 vccd1 _10355_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13117_ _16210_/Q _13120_/C _13006_/X vssd1 vssd1 vccd1 vccd1 _13117_/Y sky130_fd_sc_hd__a21oi_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14097_ _14093_/Y _14103_/A _14096_/Y _14090_/C vssd1 vssd1 vccd1 vccd1 _14099_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _13049_/B _13049_/C _13049_/A vssd1 vssd1 vccd1 vccd1 _13050_/B sky130_fd_sc_hd__a21o_1
XFILLER_112_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14999_ _15053_/A _14999_/B _15003_/B vssd1 vssd1 vccd1 vccd1 _16484_/D sky130_fd_sc_hd__nor3_1
XFILLER_47_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16738_ _16738_/A _07845_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09210_ _15569_/Q _15568_/Q _15567_/Q _09090_/X vssd1 vssd1 vccd1 vccd1 _15579_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09141_ _09141_/A _09141_/B _09141_/C vssd1 vssd1 vccd1 vccd1 _09142_/C sky130_fd_sc_hd__nand3_1
X_09072_ _09072_/A _09072_/B vssd1 vssd1 vccd1 vccd1 _09073_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08023_ _16560_/Q vssd1 vssd1 vccd1 vccd1 _11004_/A sky130_fd_sc_hd__clkinv_2
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _09744_/X _09972_/B _09973_/Y vssd1 vssd1 vccd1 vccd1 _15729_/D sky130_fd_sc_hd__o21a_1
XFILLER_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08925_ _08923_/X _08920_/A _08924_/X vssd1 vssd1 vccd1 vccd1 _08926_/B sky130_fd_sc_hd__o21ai_1
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08856_ _14858_/A vssd1 vssd1 vccd1 vccd1 _10782_/B sky130_fd_sc_hd__buf_4
XFILLER_111_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07807_ _07811_/A vssd1 vssd1 vccd1 vccd1 _07807_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08787_ _08630_/X _08780_/B _08783_/B _08786_/Y vssd1 vssd1 vccd1 vccd1 _15485_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09408_ _15620_/Q _09416_/C _09362_/X vssd1 vssd1 vccd1 vccd1 _09412_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ _10681_/B _10681_/C _10681_/A vssd1 vssd1 vccd1 vccd1 _10682_/B sky130_fd_sc_hd__a21o_1
XFILLER_139_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09339_ _09336_/A _09335_/Y _09336_/B vssd1 vssd1 vccd1 vccd1 _09339_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ _12371_/A _12350_/B _12354_/B vssd1 vssd1 vccd1 vccd1 _16099_/D sky130_fd_sc_hd__nor3_1
X_11301_ _15953_/Q _11353_/B _11301_/C vssd1 vssd1 vccd1 vccd1 _11301_/X sky130_fd_sc_hd__and3_1
X_12281_ _12276_/Y _12279_/X _12280_/Y _12274_/C vssd1 vssd1 vccd1 vccd1 _12283_/B
+ sky130_fd_sc_hd__o211ai_1
X_11232_ _11268_/C vssd1 vssd1 vccd1 vccd1 _11275_/C sky130_fd_sc_hd__clkbuf_2
X_14020_ _14035_/A _14020_/B _14020_/C vssd1 vssd1 vccd1 vccd1 _14021_/A sky130_fd_sc_hd__and3_1
X_11163_ _11163_/A _11163_/B vssd1 vssd1 vccd1 vccd1 _11164_/B sky130_fd_sc_hd__nor2_1
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10114_ _10322_/A _10114_/B vssd1 vssd1 vccd1 vccd1 _10114_/Y sky130_fd_sc_hd__nor2_1
X_15971_ _16005_/CLK _15971_/D vssd1 vssd1 vccd1 vccd1 _15971_/Q sky130_fd_sc_hd__dfxtp_1
X_11094_ _15923_/Q _11212_/B _11099_/C vssd1 vssd1 vccd1 vccd1 _11094_/Y sky130_fd_sc_hd__nand3_1
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10045_ _15746_/Q _10301_/C _10051_/C vssd1 vssd1 vccd1 vccd1 _10045_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14922_ _14922_/A vssd1 vssd1 vccd1 vccd1 _16472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14853_ _16463_/Q _14853_/B _14860_/C vssd1 vssd1 vccd1 vccd1 _14855_/C sky130_fd_sc_hd__nand3_1
XFILLER_76_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13804_ _13804_/A vssd1 vssd1 vccd1 vccd1 _16305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14784_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14909_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ _11992_/Y _11994_/X _11995_/Y _11990_/C vssd1 vssd1 vccd1 vccd1 _11998_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16523_ _16607_/CLK _16523_/D vssd1 vssd1 vccd1 vccd1 _16523_/Q sky130_fd_sc_hd__dfxtp_1
X_13735_ _13735_/A vssd1 vssd1 vccd1 vccd1 _16295_/D sky130_fd_sc_hd__clkbuf_1
X_10947_ _16559_/Q vssd1 vssd1 vccd1 vccd1 _10963_/C sky130_fd_sc_hd__inv_2
XFILLER_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16454_ input11/X _16454_/D vssd1 vssd1 vccd1 vccd1 _16454_/Q sky130_fd_sc_hd__dfxtp_1
X_13666_ _13784_/A _13666_/B _13670_/A vssd1 vssd1 vccd1 vccd1 _16286_/D sky130_fd_sc_hd__nor3_1
X_10878_ _15893_/Q _11099_/B _10878_/C vssd1 vssd1 vccd1 vccd1 _10886_/B sky130_fd_sc_hd__and3_1
X_15405_ _16125_/Q _16124_/Q _16123_/Q _15403_/X vssd1 vssd1 vccd1 vccd1 _16586_/D
+ sky130_fd_sc_hd__o31a_1
X_12617_ _12625_/A _12617_/B _12617_/C vssd1 vssd1 vccd1 vccd1 _12618_/A sky130_fd_sc_hd__and3_1
X_16385_ _16389_/CLK _16385_/D vssd1 vssd1 vccd1 vccd1 _16385_/Q sky130_fd_sc_hd__dfxtp_1
X_13597_ _13595_/A _13595_/B _13596_/X vssd1 vssd1 vccd1 vccd1 _16276_/D sky130_fd_sc_hd__a21oi_1
XFILLER_129_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15336_ _15337_/B _15337_/C _15337_/A vssd1 vssd1 vccd1 vccd1 _15338_/B sky130_fd_sc_hd__a21o_1
X_12548_ _12565_/A _12548_/B _12548_/C vssd1 vssd1 vccd1 vccd1 _12549_/A sky130_fd_sc_hd__and3_1
XFILLER_117_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15267_ _16531_/Q _15267_/B _15267_/C vssd1 vssd1 vccd1 vccd1 _15274_/B sky130_fd_sc_hd__and3_1
XANTENNA_2 _07830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12514_/A _12479_/B _12483_/A vssd1 vssd1 vccd1 vccd1 _16118_/D sky130_fd_sc_hd__nor3_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14218_ _14256_/A _14218_/B _14218_/C vssd1 vssd1 vccd1 vccd1 _14219_/A sky130_fd_sc_hd__and3_1
XFILLER_144_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15198_ _15205_/A _15198_/B _15198_/C vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__and3_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14149_ _16355_/Q _14318_/B _14154_/C vssd1 vssd1 vccd1 vccd1 _14149_/Y sky130_fd_sc_hd__nand3_1
XFILLER_140_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08710_ _08710_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _15469_/D sky130_fd_sc_hd__nor2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _09688_/A _09688_/B _09687_/Y _09689_/Y vssd1 vssd1 vccd1 vccd1 _15673_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_39_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08641_ _10016_/A vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08572_ _15232_/B vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__buf_6
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09124_ _09124_/A _09124_/B _09124_/C vssd1 vssd1 vccd1 vccd1 _09128_/A sky130_fd_sc_hd__and3_1
XFILLER_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09055_ _15549_/Q _09057_/C _09014_/X vssd1 vssd1 vccd1 vccd1 _09059_/B sky130_fd_sc_hd__a21o_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08006_ _16582_/Q vssd1 vssd1 vccd1 vccd1 _12247_/A sky130_fd_sc_hd__inv_2
XFILLER_116_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09957_ _09950_/C _09951_/C _09954_/Y _09961_/A vssd1 vssd1 vccd1 vccd1 _09961_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08908_ _08908_/A _08908_/B vssd1 vssd1 vccd1 vccd1 _08911_/A sky130_fd_sc_hd__or2_1
XFILLER_58_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09883_/Y _09886_/X _09887_/Y vssd1 vssd1 vccd1 vccd1 _15710_/D sky130_fd_sc_hd__o21a_1
XFILLER_100_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08839_ _08796_/X _08838_/A _08711_/X vssd1 vssd1 vccd1 vccd1 _08839_/Y sky130_fd_sc_hd__a21oi_1
X_16681__86 vssd1 vssd1 vccd1 vccd1 _16681__86/HI _16757_/A sky130_fd_sc_hd__conb_1
X_11850_ _11850_/A vssd1 vssd1 vccd1 vccd1 _11850_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10801_ _10801_/A _10801_/B _10801_/C vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__and3_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11781_ _11778_/Y _11787_/A _11780_/Y _11776_/C vssd1 vssd1 vccd1 vccd1 _11783_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13520_ _16267_/Q _13631_/B _13531_/C vssd1 vssd1 vccd1 vccd1 _13520_/X sky130_fd_sc_hd__and3_1
X_10732_ _10738_/A _10732_/B _10732_/C vssd1 vssd1 vccd1 vccd1 _10733_/A sky130_fd_sc_hd__and3_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13451_ _16257_/Q _13459_/C _13450_/X vssd1 vssd1 vccd1 vccd1 _13451_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10663_ _10661_/A _10661_/B _10662_/X vssd1 vssd1 vccd1 vccd1 _15855_/D sky130_fd_sc_hd__a21oi_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12402_ _16108_/Q _12456_/B _12402_/C vssd1 vssd1 vccd1 vccd1 _12411_/A sky130_fd_sc_hd__and3_1
X_16170_ _16237_/CLK _16170_/D vssd1 vssd1 vccd1 vccd1 _16170_/Q sky130_fd_sc_hd__dfxtp_1
X_13382_ _16247_/Q _13424_/C _13216_/X vssd1 vssd1 vccd1 vccd1 _13384_/B sky130_fd_sc_hd__a21oi_1
X_10594_ _10592_/Y _10593_/X _10588_/C _10589_/C vssd1 vssd1 vccd1 vccd1 _10596_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_127_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15121_ _15121_/A vssd1 vssd1 vccd1 vccd1 _15135_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12333_ _12330_/Y _12331_/X _12332_/Y _12328_/C vssd1 vssd1 vccd1 vccd1 _12335_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15052_ _15050_/Y _15045_/C _15047_/Y _15057_/A vssd1 vssd1 vccd1 vccd1 _15057_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_142_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12264_ _12260_/Y _12263_/X _12257_/C _12258_/C vssd1 vssd1 vccd1 vccd1 _12266_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_141_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14003_ _14038_/C vssd1 vssd1 vccd1 vccd1 _14044_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_135_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11215_ _11236_/A _11215_/B _11219_/B vssd1 vssd1 vccd1 vccd1 _15939_/D sky130_fd_sc_hd__nor3_1
X_12195_ _16079_/Q _12252_/B _12204_/C vssd1 vssd1 vccd1 vccd1 _12200_/A sky130_fd_sc_hd__and3_1
X_11146_ _11142_/Y _11144_/X _11145_/Y _11140_/C vssd1 vssd1 vccd1 vccd1 _11148_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_96_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15954_ _16005_/CLK _15954_/D vssd1 vssd1 vccd1 vccd1 _15954_/Q sky130_fd_sc_hd__dfxtp_1
X_11077_ _11360_/A vssd1 vssd1 vccd1 vccd1 _11309_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_110_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10028_ _15744_/Q _10057_/C _09943_/X vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__a21oi_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14905_ _14940_/C vssd1 vssd1 vccd1 vccd1 _14947_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15885_ _16570_/CLK _15885_/D vssd1 vssd1 vccd1 vccd1 _15885_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14836_ _14834_/A _14834_/B _14835_/X vssd1 vssd1 vccd1 vccd1 _16458_/D sky130_fd_sc_hd__a21oi_1
XFILLER_17_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14767_ _14765_/Y _14760_/C _14762_/Y _14772_/A vssd1 vssd1 vccd1 vccd1 _14772_/B
+ sky130_fd_sc_hd__a211oi_1
X_11979_ _16049_/Q _12204_/B _11979_/C vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__and3_1
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16506_ _16607_/CLK _16506_/D vssd1 vssd1 vccd1 vccd1 _16506_/Q sky130_fd_sc_hd__dfxtp_2
X_13718_ _13756_/A _13718_/B _13718_/C vssd1 vssd1 vccd1 vccd1 _13719_/A sky130_fd_sc_hd__and3_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14698_ _14695_/Y _14696_/X _14697_/Y _14692_/C vssd1 vssd1 vccd1 vccd1 _14700_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16437_ _16595_/CLK _16437_/D vssd1 vssd1 vccd1 vccd1 _16437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13649_ _13649_/A _13649_/B vssd1 vssd1 vccd1 vccd1 _13656_/C sky130_fd_sc_hd__nor2_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16368_ _16389_/CLK _16368_/D vssd1 vssd1 vccd1 vccd1 _16368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15319_ _15316_/Y _15317_/Y _15318_/Y vssd1 vssd1 vccd1 vccd1 _16540_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16299_ _16346_/CLK _16299_/D vssd1 vssd1 vccd1 vccd1 _16299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09811_ _09811_/A vssd1 vssd1 vccd1 vccd1 _15698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ _09737_/Y _09741_/X _09651_/X vssd1 vssd1 vccd1 vccd1 _09742_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09673_ _09674_/B _09674_/C _09674_/A vssd1 vssd1 vccd1 vccd1 _09675_/B sky130_fd_sc_hd__a21o_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08622_/A _08622_/B _08623_/X vssd1 vssd1 vccd1 vccd1 _15457_/D sky130_fd_sc_hd__a21oi_1
XFILLER_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _08555_/A vssd1 vssd1 vccd1 vccd1 _08555_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08486_ _08419_/A _08421_/X _08419_/B vssd1 vssd1 vccd1 vccd1 _08487_/B sky130_fd_sc_hd__a21bo_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ _09101_/C _09102_/C _09104_/Y _09112_/A vssd1 vssd1 vccd1 vccd1 _09112_/B
+ sky130_fd_sc_hd__a211oi_1
X_09038_ _09038_/A vssd1 vssd1 vccd1 vccd1 _09038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11000_ _11001_/B _11001_/C _10999_/X vssd1 vssd1 vccd1 vccd1 _11002_/B sky130_fd_sc_hd__o21ai_1
XFILLER_77_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ _16186_/Q _13059_/B _12952_/C vssd1 vssd1 vccd1 vccd1 _12951_/X sky130_fd_sc_hd__and3_1
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ _11900_/A _11900_/B _11901_/X vssd1 vssd1 vccd1 vccd1 _16036_/D sky130_fd_sc_hd__a21oi_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15670_ _15791_/CLK _15670_/D vssd1 vssd1 vccd1 vccd1 _15670_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12882_ _12883_/B _12883_/C _12883_/A vssd1 vssd1 vccd1 vccd1 _12884_/B sky130_fd_sc_hd__a21o_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14906_/A vssd1 vssd1 vccd1 vccd1 _14621_/X sky130_fd_sc_hd__buf_2
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _11833_/A vssd1 vssd1 vccd1 vccd1 _16026_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14550_/A _14550_/B _14551_/X vssd1 vssd1 vccd1 vccd1 _16413_/D sky130_fd_sc_hd__a21oi_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _16017_/Q _11878_/B _11764_/C vssd1 vssd1 vccd1 vccd1 _11764_/Y sky130_fd_sc_hd__nand3_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13503_/A _13503_/B _13503_/C vssd1 vssd1 vccd1 vccd1 _13504_/C sky130_fd_sc_hd__nand3_1
XFILLER_14_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10715_ _09301_/X _10708_/B _10711_/B _10714_/Y vssd1 vssd1 vccd1 vccd1 _15865_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14483_ _14481_/Y _14476_/C _14478_/Y _14488_/A vssd1 vssd1 vccd1 vccd1 _14488_/B
+ sky130_fd_sc_hd__a211oi_1
X_11695_ _11695_/A vssd1 vssd1 vccd1 vccd1 _16007_/D sky130_fd_sc_hd__clkbuf_1
X_16222_ _16261_/CLK _16222_/D vssd1 vssd1 vccd1 vccd1 _16222_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13434_ _13434_/A vssd1 vssd1 vccd1 vccd1 _16253_/D sky130_fd_sc_hd__clkbuf_1
X_10646_ _15854_/Q _10646_/B _10652_/C vssd1 vssd1 vccd1 vccd1 _10646_/Y sky130_fd_sc_hd__nand3_1
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16153_ _16555_/Q _16153_/D vssd1 vssd1 vccd1 vccd1 _16153_/Q sky130_fd_sc_hd__dfxtp_1
X_13365_ _13365_/A _13374_/B vssd1 vssd1 vccd1 vccd1 _13368_/A sky130_fd_sc_hd__or2_1
X_10577_ _15830_/Q _15829_/Q _15828_/Q _10476_/X vssd1 vssd1 vccd1 vccd1 _15840_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ _16502_/Q _15156_/B _15109_/C vssd1 vssd1 vccd1 vccd1 _15104_/Y sky130_fd_sc_hd__nand3_1
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12316_ _13443_/A vssd1 vssd1 vccd1 vccd1 _12316_/X sky130_fd_sc_hd__clkbuf_2
X_16084_ _16554_/Q _16084_/D vssd1 vssd1 vccd1 vccd1 _16084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13296_ _13296_/A vssd1 vssd1 vccd1 vccd1 _16233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15035_ _16491_/Q _15248_/B _15035_/C vssd1 vssd1 vccd1 vccd1 _15035_/Y sky130_fd_sc_hd__nand3_1
X_12247_ _12247_/A vssd1 vssd1 vccd1 vccd1 _12263_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _16077_/Q _12179_/C _12007_/X vssd1 vssd1 vccd1 vccd1 _12180_/A sky130_fd_sc_hd__a21oi_1
X_11129_ _11126_/Y _11128_/X _11123_/C _11124_/C vssd1 vssd1 vccd1 vccd1 _11131_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15937_ _16005_/CLK _15937_/D vssd1 vssd1 vccd1 vccd1 _15937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15868_ _16570_/CLK _15868_/D vssd1 vssd1 vccd1 vccd1 _15868_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14819_ _14819_/A _14819_/B _14819_/C vssd1 vssd1 vccd1 vccd1 _14820_/A sky130_fd_sc_hd__and3_1
X_15799_ _15812_/CLK _15799_/D vssd1 vssd1 vccd1 vccd1 _15799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08340_ _08138_/A _08340_/B vssd1 vssd1 vccd1 vccd1 _08340_/X sky130_fd_sc_hd__and2b_1
XFILLER_149_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08271_ _08090_/A _08090_/B _08270_/Y vssd1 vssd1 vccd1 vccd1 _08273_/B sky130_fd_sc_hd__o21a_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07986_ _13886_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07987_/B sky130_fd_sc_hd__nand2_1
X_09725_ _09953_/A vssd1 vssd1 vccd1 vccd1 _09841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09656_ _09656_/A _09656_/B vssd1 vssd1 vccd1 vccd1 _09656_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16651__56 vssd1 vssd1 vccd1 vccd1 _16651__56/HI _16727_/A sky130_fd_sc_hd__conb_1
X_08607_ _09998_/B vssd1 vssd1 vccd1 vccd1 _10743_/B sky130_fd_sc_hd__buf_2
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09587_ _09587_/A _09587_/B _09587_/C vssd1 vssd1 vccd1 vccd1 _09588_/C sky130_fd_sc_hd__nand3_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08538_/A _08499_/B vssd1 vssd1 vccd1 vccd1 _08540_/A sky130_fd_sc_hd__or2b_1
X_08469_ _08469_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08469_/Y sky130_fd_sc_hd__nor2_1
X_10500_ _15828_/Q _10509_/C _10393_/X vssd1 vssd1 vccd1 vccd1 _10500_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11480_ _15977_/Q _11594_/B _11480_/C vssd1 vssd1 vccd1 vccd1 _11480_/Y sky130_fd_sc_hd__nand3_1
XFILLER_137_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10431_ _10740_/A vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13150_ _13151_/B _13151_/C _12982_/X vssd1 vssd1 vccd1 vccd1 _13152_/B sky130_fd_sc_hd__o21ai_1
X_10362_ _15803_/Q _10463_/B _10362_/C vssd1 vssd1 vccd1 vccd1 _10363_/B sky130_fd_sc_hd__and3_1
XFILLER_136_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12101_ _12098_/Y _12099_/X _12100_/Y _12096_/C vssd1 vssd1 vccd1 vccd1 _12103_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10293_ _15791_/Q _10294_/B _10243_/X vssd1 vssd1 vccd1 vccd1 _10293_/Y sky130_fd_sc_hd__a21oi_1
X_13081_ _16205_/Q _13082_/C _12857_/X vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__a21oi_1
XFILLER_124_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12032_ _12033_/B _12033_/C _12033_/A vssd1 vssd1 vccd1 vccd1 _12034_/B sky130_fd_sc_hd__a21o_1
XFILLER_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13983_ _13980_/Y _13991_/A _13982_/Y _13977_/C vssd1 vssd1 vccd1 vccd1 _13985_/B
+ sky130_fd_sc_hd__o211a_1
X_15722_ _15812_/CLK _15722_/D vssd1 vssd1 vccd1 vccd1 _15722_/Q sky130_fd_sc_hd__dfxtp_1
X_12934_ _16183_/Q _12975_/C _12933_/X vssd1 vssd1 vccd1 vccd1 _12936_/B sky130_fd_sc_hd__a21oi_1
XFILLER_18_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15653_ _15791_/CLK _15653_/D vssd1 vssd1 vccd1 vccd1 _15653_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12865_ _12863_/A _12863_/B _12864_/X vssd1 vssd1 vccd1 vccd1 _16172_/D sky130_fd_sc_hd__a21oi_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14604_ _14604_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14606_/A sky130_fd_sc_hd__or2_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _11810_/C _11811_/C _11813_/Y _11814_/X vssd1 vssd1 vccd1 vccd1 _11817_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _16551_/CLK _15584_/D vssd1 vssd1 vccd1 vccd1 _15584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12796_/A _12796_/B _12800_/B vssd1 vssd1 vccd1 vccd1 _16163_/D sky130_fd_sc_hd__nor3_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14535_/A _14535_/B _14535_/C vssd1 vssd1 vccd1 vccd1 _14536_/A sky130_fd_sc_hd__and3_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11805_/A _11747_/B _11752_/A vssd1 vssd1 vccd1 vccd1 _16014_/D sky130_fd_sc_hd__nor3_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14466_ _16401_/Q _14697_/B _14466_/C vssd1 vssd1 vccd1 vccd1 _14466_/Y sky130_fd_sc_hd__nand3_1
X_11678_ _11679_/B _11679_/C _11567_/X vssd1 vssd1 vccd1 vccd1 _11680_/B sky130_fd_sc_hd__o21ai_1
X_16205_ _16237_/CLK _16205_/D vssd1 vssd1 vccd1 vccd1 _16205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ _16251_/Q _13474_/B _13424_/C vssd1 vssd1 vccd1 vccd1 _13417_/Y sky130_fd_sc_hd__nand3_1
X_10629_ _15852_/Q _10658_/C _10426_/X vssd1 vssd1 vccd1 vccd1 _10631_/B sky130_fd_sc_hd__a21oi_1
X_14397_ _16391_/Q _14506_/B _14406_/C vssd1 vssd1 vccd1 vccd1 _14402_/A sky130_fd_sc_hd__and3_1
X_16136_ _16261_/CLK _16136_/D vssd1 vssd1 vccd1 vccd1 _16136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13348_ _13348_/A vssd1 vssd1 vccd1 vccd1 _16241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16067_ _16118_/CLK _16067_/D vssd1 vssd1 vccd1 vccd1 _16067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13279_ _13279_/A _13279_/B _13279_/C vssd1 vssd1 vccd1 vccd1 _13280_/C sky130_fd_sc_hd__nand3_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15018_ _16489_/Q _15074_/B _15027_/C vssd1 vssd1 vccd1 vccd1 _15023_/A sky130_fd_sc_hd__and3_1
XFILLER_111_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07840_ _07842_/A vssd1 vssd1 vccd1 vccd1 _07840_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07771_ _07774_/A vssd1 vssd1 vccd1 vccd1 _07771_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09510_ _09595_/A _09510_/B _09513_/B vssd1 vssd1 vccd1 vccd1 _15636_/D sky130_fd_sc_hd__nor3_1
XFILLER_37_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _09394_/X _09436_/B _09351_/X vssd1 vssd1 vccd1 vccd1 _09443_/A sky130_fd_sc_hd__a21oi_1
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09372_ _09370_/Y _09377_/A _09366_/C _09367_/C vssd1 vssd1 vccd1 vccd1 _09374_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08323_ _08323_/A _08196_/A vssd1 vssd1 vccd1 vccd1 _08323_/X sky130_fd_sc_hd__or2b_1
X_08254_ _08254_/A vssd1 vssd1 vccd1 vccd1 _08978_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_138_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08185_ _08186_/A _08186_/B _08186_/C vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__a21o_1
XFILLER_118_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07969_ _10767_/A _08191_/B vssd1 vssd1 vccd1 vccd1 _07970_/B sky130_fd_sc_hd__xnor2_2
X_09708_ _09617_/X _09706_/X _09701_/B _09707_/X vssd1 vssd1 vccd1 vccd1 _09709_/B
+ sky130_fd_sc_hd__a31o_1
X_10980_ _10978_/Y _10973_/C _10975_/Y _10976_/X vssd1 vssd1 vccd1 vccd1 _10981_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09639_ _09718_/A _09639_/B _09642_/B vssd1 vssd1 vccd1 vccd1 _15663_/D sky130_fd_sc_hd__nor3_1
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12650_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__buf_2
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11601_ _15994_/Q _11773_/B _11607_/C vssd1 vssd1 vccd1 vccd1 _11601_/Y sky130_fd_sc_hd__nand3_1
XFILLER_24_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12581_ _12581_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12586_/C sky130_fd_sc_hd__nor2_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14320_ _14318_/Y _14314_/C _14316_/Y _14325_/A vssd1 vssd1 vccd1 vccd1 _14325_/B
+ sky130_fd_sc_hd__a211oi_1
X_11532_ _11547_/A _11532_/B _11532_/C vssd1 vssd1 vccd1 vccd1 _11533_/A sky130_fd_sc_hd__and3_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ _14814_/A vssd1 vssd1 vccd1 vccd1 _14472_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11463_ _12029_/A vssd1 vssd1 vccd1 vccd1 _11463_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ _13202_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _13209_/C sky130_fd_sc_hd__nor2_1
XFILLER_139_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10414_ _10414_/A vssd1 vssd1 vccd1 vccd1 _10414_/X sky130_fd_sc_hd__clkbuf_2
X_14182_ _14197_/A _14182_/B _14182_/C vssd1 vssd1 vccd1 vccd1 _14183_/A sky130_fd_sc_hd__and3_1
X_11394_ _13085_/A vssd1 vssd1 vccd1 vccd1 _14220_/A sky130_fd_sc_hd__buf_6
XFILLER_136_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13133_ _13979_/A vssd1 vssd1 vccd1 vccd1 _13133_/X sky130_fd_sc_hd__buf_2
XFILLER_124_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ _10399_/A _10345_/B _10345_/C vssd1 vssd1 vccd1 vccd1 _10346_/A sky130_fd_sc_hd__and3_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _13062_/Y _13056_/C _13058_/Y _13059_/X vssd1 vssd1 vccd1 vccd1 _13065_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_140_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10276_ _10276_/A vssd1 vssd1 vccd1 vccd1 _10276_/X sky130_fd_sc_hd__clkbuf_2
X_12015_ _12013_/A _12013_/B _12014_/X vssd1 vssd1 vccd1 vccd1 _16052_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16754_ _16754_/A _07772_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
X_13966_ _16329_/Q _14135_/B _13966_/C vssd1 vssd1 vccd1 vccd1 _13966_/Y sky130_fd_sc_hd__nand3_1
XFILLER_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15705_ _15791_/CLK _15705_/D vssd1 vssd1 vccd1 vccd1 _15705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12917_ _12917_/A _12925_/B vssd1 vssd1 vccd1 vccd1 _12919_/A sky130_fd_sc_hd__or2_1
X_13897_ _13918_/A _13897_/B _13897_/C vssd1 vssd1 vccd1 vccd1 _13898_/A sky130_fd_sc_hd__and3_1
X_15636_ _15791_/CLK _15636_/D vssd1 vssd1 vccd1 vccd1 _15636_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ _12848_/A vssd1 vssd1 vccd1 vccd1 _16170_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15567_ _16551_/CLK _15567_/D vssd1 vssd1 vccd1 vccd1 _15567_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _12775_/Y _12776_/X _12778_/Y _12773_/C vssd1 vssd1 vccd1 vccd1 _12781_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14518_ _14511_/C _14512_/C _14514_/Y _14516_/X vssd1 vssd1 vccd1 vccd1 _14519_/C
+ sky130_fd_sc_hd__a211o_1
X_15498_ _16570_/CLK _15498_/D vssd1 vssd1 vccd1 vccd1 _15498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14449_ _16399_/Q _14506_/B _14458_/C vssd1 vssd1 vccd1 vccd1 _14454_/A sky130_fd_sc_hd__and3_1
XFILLER_128_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16119_ _16554_/Q _16119_/D vssd1 vssd1 vccd1 vccd1 _16119_/Q sky130_fd_sc_hd__dfxtp_1
X_09990_ _10340_/A vssd1 vssd1 vccd1 vccd1 _10082_/A sky130_fd_sc_hd__buf_2
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08941_ _08941_/A vssd1 vssd1 vccd1 vccd1 _15518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _09076_/A vssd1 vssd1 vccd1 vccd1 _08872_/X sky130_fd_sc_hd__buf_2
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07823_ _07824_/A vssd1 vssd1 vccd1 vccd1 _07823_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16621__26 vssd1 vssd1 vccd1 vccd1 _16621__26/HI _16687_/A sky130_fd_sc_hd__conb_1
X_09424_ _09698_/A vssd1 vssd1 vccd1 vccd1 _09424_/X sky130_fd_sc_hd__buf_2
XFILLER_52_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ _15740_/Q _15739_/Q _15738_/Q _09314_/X vssd1 vssd1 vccd1 vccd1 _15606_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ _08306_/A _08306_/B vssd1 vssd1 vccd1 vccd1 _15293_/C sky130_fd_sc_hd__xor2_2
X_09286_ _15596_/Q _09472_/B _09286_/C vssd1 vssd1 vccd1 vccd1 _09286_/X sky130_fd_sc_hd__and3_1
X_08237_ _08237_/A _08237_/B vssd1 vssd1 vccd1 vccd1 _08238_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08168_ _13551_/A _07943_/B _08167_/Y vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__o21a_1
XFILLER_119_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08099_ _15570_/Q _08292_/B vssd1 vssd1 vccd1 vccd1 _08100_/B sky130_fd_sc_hd__xnor2_2
X_10130_ _10145_/A _10130_/B _10130_/C vssd1 vssd1 vccd1 vccd1 _10131_/A sky130_fd_sc_hd__and3_1
XFILLER_133_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10061_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10062_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13820_ _13927_/A _13820_/B _13824_/B vssd1 vssd1 vccd1 vccd1 _16307_/D sky130_fd_sc_hd__nor3_1
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ _16299_/Q _13759_/C _13750_/X vssd1 vssd1 vccd1 vccd1 _13751_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10963_ _15905_/Q _11070_/B _10963_/C vssd1 vssd1 vccd1 vccd1 _10963_/X sky130_fd_sc_hd__and3_1
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12702_ _12736_/A _12702_/B _12702_/C vssd1 vssd1 vccd1 vccd1 _12703_/A sky130_fd_sc_hd__and3_1
X_16470_ input11/X _16470_/D vssd1 vssd1 vccd1 vccd1 _16470_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13682_ _13682_/A vssd1 vssd1 vccd1 vccd1 _13906_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10894_ _15232_/B vssd1 vssd1 vccd1 vccd1 _11118_/B sky130_fd_sc_hd__buf_2
XFILLER_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15421_ _16229_/Q _16228_/Q _16227_/Q _15416_/X vssd1 vssd1 vccd1 vccd1 _16599_/D
+ sky130_fd_sc_hd__o31a_1
X_12633_ _16141_/Q _12634_/C _12575_/X vssd1 vssd1 vccd1 vccd1 _12635_/A sky130_fd_sc_hd__a21oi_1
XFILLER_43_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15352_ _15347_/B _15350_/B _09117_/X vssd1 vssd1 vccd1 vccd1 _15358_/C sky130_fd_sc_hd__o21a_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12564_ _12562_/Y _12557_/C _12559_/Y _12561_/X vssd1 vssd1 vccd1 vccd1 _12565_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303_ _16377_/Q _14414_/B _14303_/C vssd1 vssd1 vccd1 vccd1 _14303_/Y sky130_fd_sc_hd__nand3_1
X_11515_ _11551_/C vssd1 vssd1 vccd1 vccd1 _11560_/C sky130_fd_sc_hd__clkbuf_2
X_15283_ _15333_/A _15283_/B _15283_/C vssd1 vssd1 vccd1 vccd1 _16535_/D sky130_fd_sc_hd__nor3_1
X_12495_ _16121_/Q _12726_/B _12495_/C vssd1 vssd1 vccd1 vccd1 _12495_/Y sky130_fd_sc_hd__nand3_1
X_14234_ _14234_/A vssd1 vssd1 vccd1 vccd1 _16367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11446_ _11446_/A _11446_/B vssd1 vssd1 vccd1 vccd1 _11447_/B sky130_fd_sc_hd__nor2_1
XFILLER_125_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14165_ _16616_/Q vssd1 vssd1 vccd1 vccd1 _14179_/C sky130_fd_sc_hd__clkinv_2
X_11377_ _11373_/Y _11383_/A _11376_/Y _11371_/C vssd1 vssd1 vccd1 vccd1 _11379_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ _13116_/A vssd1 vssd1 vccd1 vccd1 _16208_/D sky130_fd_sc_hd__clkbuf_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _10332_/C vssd1 vssd1 vccd1 vccd1 _10342_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14096_ _16347_/Q _14318_/B _14101_/C vssd1 vssd1 vccd1 vccd1 _14096_/Y sky130_fd_sc_hd__nand3_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _16200_/Q _13164_/B _13053_/C vssd1 vssd1 vccd1 vccd1 _13049_/C sky130_fd_sc_hd__nand3_1
XFILLER_140_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10259_ _10259_/A vssd1 vssd1 vccd1 vccd1 _15781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14998_ _14996_/Y _14992_/C _14994_/Y _15003_/A vssd1 vssd1 vccd1 vccd1 _15003_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16737_ _16737_/A _07844_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13949_ _14063_/A _13949_/B _13953_/A vssd1 vssd1 vccd1 vccd1 _16326_/D sky130_fd_sc_hd__nor3_1
XFILLER_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ _15812_/CLK _15619_/D vssd1 vssd1 vccd1 vccd1 _15619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16599_ _16607_/CLK _16599_/D vssd1 vssd1 vccd1 vccd1 _16599_/Q sky130_fd_sc_hd__dfxtp_1
X_09140_ _09141_/B _09141_/C _09141_/A vssd1 vssd1 vccd1 vccd1 _09142_/B sky130_fd_sc_hd__a21o_1
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09071_ _09071_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09073_/A sky130_fd_sc_hd__or2_1
X_08022_ _10076_/C _08022_/B vssd1 vssd1 vccd1 vccd1 _08096_/A sky130_fd_sc_hd__xnor2_2
XFILLER_128_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09973_ _10017_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _09973_/Y sky130_fd_sc_hd__nor2_1
X_08924_ _15338_/A vssd1 vssd1 vccd1 vccd1 _08924_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08855_ input2/X vssd1 vssd1 vccd1 vccd1 _14858_/A sky130_fd_sc_hd__buf_2
XFILLER_85_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07806_ _07806_/A vssd1 vssd1 vccd1 vccd1 _07811_/A sky130_fd_sc_hd__clkbuf_4
X_08786_ _08916_/A _08791_/C vssd1 vssd1 vccd1 vccd1 _08786_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09407_ _09812_/A vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09338_ _09336_/A _09336_/B _09335_/Y _09337_/Y vssd1 vssd1 vccd1 vccd1 _15601_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_138_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ _09261_/C _09262_/C _09265_/Y _09276_/A vssd1 vssd1 vccd1 vccd1 _09276_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11300_ _15953_/Q _11309_/C _11188_/X vssd1 vssd1 vccd1 vccd1 _11300_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12280_ _16090_/Q _12340_/B _12287_/C vssd1 vssd1 vccd1 vccd1 _12280_/Y sky130_fd_sc_hd__nand3_1
X_11231_ _11253_/C vssd1 vssd1 vccd1 vccd1 _11268_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11162_ _11162_/A _11169_/B vssd1 vssd1 vccd1 vccd1 _11164_/A sky130_fd_sc_hd__or2_1
XFILLER_134_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10113_ _10107_/B _10110_/B _09125_/A vssd1 vssd1 vccd1 vccd1 _10114_/B sky130_fd_sc_hd__o21a_1
XFILLER_121_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15970_ _16005_/CLK _15970_/D vssd1 vssd1 vccd1 vccd1 _15970_/Q sky130_fd_sc_hd__dfxtp_1
X_11093_ _15924_/Q _11322_/B _11093_/C vssd1 vssd1 vccd1 vccd1 _11101_/A sky130_fd_sc_hd__and3_1
XFILLER_96_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10044_ _15747_/Q _10300_/C _10051_/C vssd1 vssd1 vccd1 vccd1 _10044_/X sky130_fd_sc_hd__and3_1
X_14921_ _14936_/A _14921_/B _14921_/C vssd1 vssd1 vccd1 vccd1 _14922_/A sky130_fd_sc_hd__and3_1
X_14852_ _16463_/Q _14860_/C _14851_/X vssd1 vssd1 vccd1 vccd1 _14855_/B sky130_fd_sc_hd__a21o_1
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13803_ _13811_/A _13803_/B _13803_/C vssd1 vssd1 vccd1 vccd1 _13804_/A sky130_fd_sc_hd__and3_1
X_14783_ _16441_/Q _16440_/Q _16439_/Q _14615_/X vssd1 vssd1 vccd1 vccd1 _16451_/D
+ sky130_fd_sc_hd__o31a_1
X_11995_ _16050_/Q _12053_/B _12002_/C vssd1 vssd1 vccd1 vccd1 _11995_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13734_ _13756_/A _13734_/B _13734_/C vssd1 vssd1 vccd1 vccd1 _13735_/A sky130_fd_sc_hd__and3_1
X_16522_ _16595_/CLK _16522_/D vssd1 vssd1 vccd1 vccd1 _16522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10946_ _10946_/A vssd1 vssd1 vccd1 vccd1 _15901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13665_ _16287_/Q _13665_/B _13676_/C vssd1 vssd1 vccd1 vccd1 _13670_/A sky130_fd_sc_hd__and3_1
X_16453_ input11/X _16453_/D vssd1 vssd1 vccd1 vccd1 _16453_/Q sky130_fd_sc_hd__dfxtp_1
X_10877_ _12009_/A vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12616_ _12614_/Y _12610_/C _12612_/Y _12613_/X vssd1 vssd1 vccd1 vccd1 _12617_/C
+ sky130_fd_sc_hd__a211o_1
X_15404_ _16117_/Q _16116_/Q _16115_/Q _15403_/X vssd1 vssd1 vccd1 vccd1 _16585_/D
+ sky130_fd_sc_hd__o31a_1
X_16384_ _16389_/CLK _16384_/D vssd1 vssd1 vccd1 vccd1 _16384_/Q sky130_fd_sc_hd__dfxtp_1
X_13596_ _13596_/A _13600_/C vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__or2_1
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ _16549_/Q _15335_/B _15335_/C vssd1 vssd1 vccd1 vccd1 _15337_/C sky130_fd_sc_hd__nand3_1
XFILLER_61_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12547_ _12540_/C _12541_/C _12543_/Y _12545_/X vssd1 vssd1 vccd1 vccd1 _12548_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15266_ _16531_/Q _15267_/C _10812_/B vssd1 vssd1 vccd1 vccd1 _15268_/A sky130_fd_sc_hd__a21oi_1
X_12478_ _16119_/Q _12535_/B _12487_/C vssd1 vssd1 vccd1 vccd1 _12483_/A sky130_fd_sc_hd__and3_1
XANTENNA_3 _07842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14217_ _14276_/A _14217_/B _14217_/C vssd1 vssd1 vccd1 vccd1 _14218_/C sky130_fd_sc_hd__or3_1
X_11429_ _11425_/Y _11427_/X _11428_/Y _11423_/C vssd1 vssd1 vccd1 vccd1 _11431_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15197_ _15195_/Y _15191_/C _15193_/Y _15194_/X vssd1 vssd1 vccd1 vccd1 _15198_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_99_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14148_ _16356_/Q _14148_/B _14148_/C vssd1 vssd1 vccd1 vccd1 _14156_/A sky130_fd_sc_hd__and3_1
XFILLER_125_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14079_ _16345_/Q _14135_/B _14079_/C vssd1 vssd1 vccd1 vccd1 _14079_/Y sky130_fd_sc_hd__nand3_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08640_ _09699_/A vssd1 vssd1 vccd1 vccd1 _10016_/A sky130_fd_sc_hd__buf_2
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08571_ input9/X vssd1 vssd1 vccd1 vccd1 _15232_/B sky130_fd_sc_hd__clkbuf_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09123_ _09123_/A _09123_/B vssd1 vssd1 vccd1 vccd1 _15558_/D sky130_fd_sc_hd__nor2_1
X_09054_ _09054_/A _09054_/B _09059_/A vssd1 vssd1 vccd1 vccd1 _15544_/D sky130_fd_sc_hd__nor3_1
X_08005_ _16558_/Q vssd1 vssd1 vccd1 vccd1 _10889_/A sky130_fd_sc_hd__inv_2
XFILLER_150_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09956_ _09954_/Y _09961_/A _09950_/C _09951_/C vssd1 vssd1 vccd1 vccd1 _09958_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08907_ _15515_/Q _08991_/B _08907_/C vssd1 vssd1 vccd1 vccd1 _08908_/B sky130_fd_sc_hd__and3_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09883_/Y _09886_/X _09750_/X vssd1 vssd1 vccd1 vccd1 _09887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08838_ _08838_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _15496_/D sky130_fd_sc_hd__nor2_1
XFILLER_73_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08769_ _08940_/A _08769_/B _08769_/C vssd1 vssd1 vccd1 vccd1 _08770_/A sky130_fd_sc_hd__and3_1
XFILLER_72_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10800_ _10798_/Y _10794_/C _10796_/Y _10797_/X vssd1 vssd1 vccd1 vccd1 _10801_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11780_ _16019_/Q _11780_/B _11785_/C vssd1 vssd1 vccd1 vccd1 _11780_/Y sky130_fd_sc_hd__nand3_1
XFILLER_26_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731_ _10731_/A _10731_/B _10731_/C vssd1 vssd1 vccd1 vccd1 _10732_/C sky130_fd_sc_hd__nand3_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13450_ _14015_/A vssd1 vssd1 vccd1 vccd1 _13450_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10662_ _10759_/A _10662_/B vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__or2_1
XFILLER_139_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _16108_/Q _12409_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12401_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13381_ _13416_/C vssd1 vssd1 vccd1 vccd1 _13424_/C sky130_fd_sc_hd__clkbuf_2
X_10593_ _15845_/Q _10735_/B _10593_/C vssd1 vssd1 vccd1 vccd1 _10593_/X sky130_fd_sc_hd__and3_1
X_15120_ _16495_/Q _16494_/Q _16493_/Q _14900_/X vssd1 vssd1 vccd1 vccd1 _16505_/D
+ sky130_fd_sc_hd__o31a_1
X_12332_ _16097_/Q _12443_/B _12332_/C vssd1 vssd1 vccd1 vccd1 _12332_/Y sky130_fd_sc_hd__nand3_1
XFILLER_126_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _15047_/Y _15057_/A _15050_/Y _15045_/C vssd1 vssd1 vccd1 vccd1 _15053_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ _16089_/Q _12487_/B _12263_/C vssd1 vssd1 vccd1 vccd1 _12263_/X sky130_fd_sc_hd__and3_1
X_14002_ _14024_/C vssd1 vssd1 vccd1 vccd1 _14038_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11214_ _11212_/Y _11208_/C _11210_/Y _11219_/A vssd1 vssd1 vccd1 vccd1 _11219_/B
+ sky130_fd_sc_hd__a211oi_1
X_12194_ _16079_/Q _12232_/C _12081_/X vssd1 vssd1 vccd1 vccd1 _12196_/B sky130_fd_sc_hd__a21oi_1
X_11145_ _15930_/Q _11205_/B _11152_/C vssd1 vssd1 vccd1 vccd1 _11145_/Y sky130_fd_sc_hd__nand3_1
XFILLER_110_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16657__62 vssd1 vssd1 vccd1 vccd1 _16657__62/HI _16733_/A sky130_fd_sc_hd__conb_1
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15953_ _15365_/A _15953_/D vssd1 vssd1 vccd1 vccd1 _15953_/Q sky130_fd_sc_hd__dfxtp_1
X_11076_ _15922_/Q _11076_/B _11078_/C vssd1 vssd1 vccd1 vccd1 _11076_/X sky130_fd_sc_hd__and3_1
XFILLER_110_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10027_ _10051_/C vssd1 vssd1 vccd1 vccd1 _10057_/C sky130_fd_sc_hd__clkbuf_2
X_14904_ _14925_/C vssd1 vssd1 vccd1 vccd1 _14940_/C sky130_fd_sc_hd__clkbuf_2
X_15884_ _16553_/Q _15884_/D vssd1 vssd1 vccd1 vccd1 _15884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14835_ _15005_/A _14839_/C vssd1 vssd1 vccd1 vccd1 _14835_/X sky130_fd_sc_hd__or2_1
XFILLER_17_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11978_ _11978_/A vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14766_ _14762_/Y _14772_/A _14765_/Y _14760_/C vssd1 vssd1 vccd1 vccd1 _14768_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _16607_/CLK _16505_/D vssd1 vssd1 vccd1 vccd1 _16505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10929_ _15899_/Q _10929_/B _10934_/C vssd1 vssd1 vccd1 vccd1 _10929_/Y sky130_fd_sc_hd__nand3_1
X_13717_ _13717_/A _13717_/B _13717_/C vssd1 vssd1 vccd1 vccd1 _13718_/C sky130_fd_sc_hd__or3_1
X_14697_ _16437_/Q _14697_/B _14697_/C vssd1 vssd1 vccd1 vccd1 _14697_/Y sky130_fd_sc_hd__nand3_1
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16436_ _16595_/CLK _16436_/D vssd1 vssd1 vccd1 vccd1 _16436_/Q sky130_fd_sc_hd__dfxtp_1
X_13648_ _14210_/A vssd1 vssd1 vccd1 vccd1 _13879_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16367_ _16389_/CLK _16367_/D vssd1 vssd1 vccd1 vccd1 _16367_/Q sky130_fd_sc_hd__dfxtp_1
X_13579_ _16275_/Q _13631_/B _13586_/C vssd1 vssd1 vccd1 vccd1 _13579_/X sky130_fd_sc_hd__and3_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15318_ _15316_/Y _15317_/Y _10716_/X vssd1 vssd1 vccd1 vccd1 _15318_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16298_ _16533_/Q _16298_/D vssd1 vssd1 vccd1 vccd1 _16298_/Q sky130_fd_sc_hd__dfxtp_1
X_15249_ _15246_/Y _15247_/X _15248_/Y _15244_/C vssd1 vssd1 vccd1 vccd1 _15251_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_99_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09810_ _09810_/A _09810_/B _09810_/C vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__and3_1
XFILLER_141_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _09739_/X _09741_/B vssd1 vssd1 vccd1 vccd1 _09741_/X sky130_fd_sc_hd__and2b_1
XFILLER_140_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09672_ _15674_/Q _09867_/B _09679_/C vssd1 vssd1 vccd1 vccd1 _09674_/C sky130_fd_sc_hd__nand3_1
XFILLER_55_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08623_ _15207_/A _08623_/B vssd1 vssd1 vccd1 vccd1 _08623_/X sky130_fd_sc_hd__or2_1
XFILLER_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _08554_/A vssd1 vssd1 vccd1 vccd1 _15366_/B sky130_fd_sc_hd__buf_6
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08485_ _08485_/A _08485_/B vssd1 vssd1 vccd1 vccd1 _08487_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09106_ _09104_/Y _09112_/A _09101_/C _09102_/C vssd1 vssd1 vccd1 vccd1 _09108_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09037_ _09037_/A _09042_/C vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__and2_1
XFILLER_136_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09939_ _15713_/Q _15712_/Q _15711_/Q _09756_/X vssd1 vssd1 vccd1 vccd1 _15723_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12950_ _16186_/Q _12952_/C _12723_/X vssd1 vssd1 vccd1 vccd1 _12950_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11901_ _11901_/A _11905_/C vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__or2_1
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12881_ _16176_/Q _12881_/B _12889_/C vssd1 vssd1 vccd1 vccd1 _12883_/C sky130_fd_sc_hd__nand3_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _11832_/A _11832_/B _11832_/C vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__and3_1
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14620_ _14655_/C vssd1 vssd1 vccd1 vccd1 _14662_/C sky130_fd_sc_hd__clkbuf_2
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14720_/A _14555_/C vssd1 vssd1 vccd1 vccd1 _14551_/X sky130_fd_sc_hd__or2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11763_ _16018_/Q _11928_/B _11764_/C vssd1 vssd1 vccd1 vccd1 _11763_/X sky130_fd_sc_hd__and3_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13503_/B _13503_/C _13503_/A vssd1 vssd1 vccd1 vccd1 _13504_/B sky130_fd_sc_hd__a21o_1
X_10714_ _15353_/A _10714_/B vssd1 vssd1 vccd1 vccd1 _10714_/Y sky130_fd_sc_hd__nor2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14478_/Y _14488_/A _14481_/Y _14476_/C vssd1 vssd1 vccd1 vccd1 _14484_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11694_ _11717_/A _11694_/B _11694_/C vssd1 vssd1 vccd1 vccd1 _11695_/A sky130_fd_sc_hd__and3_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13433_ _13470_/A _13433_/B _13433_/C vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__and3_1
X_16221_ _16237_/CLK _16221_/D vssd1 vssd1 vccd1 vccd1 _16221_/Q sky130_fd_sc_hd__dfxtp_1
X_10645_ _15855_/Q _10691_/B _10652_/C vssd1 vssd1 vccd1 vccd1 _10645_/X sky130_fd_sc_hd__and3_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16152_ _16261_/CLK _16152_/D vssd1 vssd1 vccd1 vccd1 _16152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13364_ _16245_/Q _13364_/B _13364_/C vssd1 vssd1 vccd1 vccd1 _13374_/B sky130_fd_sc_hd__and3_1
X_10576_ _10526_/X _10573_/B _10575_/Y vssd1 vssd1 vccd1 vccd1 _15839_/D sky130_fd_sc_hd__o21a_1
X_12315_ input10/X vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__buf_4
X_15103_ _16503_/Q _15261_/B _15103_/C vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__and3_1
X_16083_ _16118_/CLK _16083_/D vssd1 vssd1 vccd1 vccd1 _16083_/Q sky130_fd_sc_hd__dfxtp_1
X_13295_ _13302_/A _13295_/B _13295_/C vssd1 vssd1 vccd1 vccd1 _13296_/A sky130_fd_sc_hd__and3_1
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15034_ _15034_/A vssd1 vssd1 vccd1 vccd1 _15248_/B sky130_fd_sc_hd__buf_2
X_12246_ _12683_/A vssd1 vssd1 vccd1 vccd1 _12371_/A sky130_fd_sc_hd__buf_2
XFILLER_142_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12177_ _12230_/A _12177_/B _12181_/B vssd1 vssd1 vccd1 vccd1 _16075_/D sky130_fd_sc_hd__nor3_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11128_ _15929_/Q _11353_/B _11128_/C vssd1 vssd1 vccd1 vccd1 _11128_/X sky130_fd_sc_hd__and3_1
XFILLER_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15936_ _16005_/CLK _15936_/D vssd1 vssd1 vccd1 vccd1 _15936_/Q sky130_fd_sc_hd__dfxtp_1
X_11059_ _11093_/C vssd1 vssd1 vccd1 vccd1 _11099_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15867_ _16595_/CLK _15867_/D vssd1 vssd1 vccd1 vccd1 _15867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14818_ _14816_/Y _14811_/C _14813_/Y _14815_/X vssd1 vssd1 vccd1 vccd1 _14819_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15798_ _16595_/CLK _15798_/D vssd1 vssd1 vccd1 vccd1 _15798_/Q sky130_fd_sc_hd__dfxtp_1
X_14749_ _15034_/A vssd1 vssd1 vccd1 vccd1 _14982_/B sky130_fd_sc_hd__buf_2
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08270_ _16592_/Q _08270_/B vssd1 vssd1 vccd1 vccd1 _08270_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16419_ _16595_/CLK _16419_/D vssd1 vssd1 vccd1 vccd1 _16419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07985_ _13886_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _08186_/B sky130_fd_sc_hd__or2_1
XFILLER_86_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09724_ _09724_/A vssd1 vssd1 vccd1 vccd1 _15680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09655_ _09655_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09656_/B sky130_fd_sc_hd__and2_1
XFILLER_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08606_ _09815_/A vssd1 vssd1 vccd1 vccd1 _09998_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09586_ _09587_/B _09587_/C _09587_/A vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__a21o_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08537_/A _08537_/B vssd1 vssd1 vccd1 vccd1 _08540_/C sky130_fd_sc_hd__nand2_1
XFILLER_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08468_ _08496_/A _08496_/B vssd1 vssd1 vccd1 vccd1 _08512_/A sky130_fd_sc_hd__xnor2_4
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08399_ _08399_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08469_/A sky130_fd_sc_hd__xnor2_4
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10430_ _10430_/A vssd1 vssd1 vccd1 vccd1 _10740_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10361_ _15803_/Q _10362_/C _10360_/X vssd1 vssd1 vccd1 vccd1 _10363_/A sky130_fd_sc_hd__a21oi_1
XFILLER_128_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12100_ _16065_/Q _12160_/B _12100_/C vssd1 vssd1 vccd1 vccd1 _12100_/Y sky130_fd_sc_hd__nand3_1
XFILLER_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ _13080_/A _13080_/B _13084_/B vssd1 vssd1 vccd1 vccd1 _16203_/D sky130_fd_sc_hd__nor3_1
XFILLER_124_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10292_ _10292_/A vssd1 vssd1 vccd1 vccd1 _15788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _16056_/Q _12031_/B _12038_/C vssd1 vssd1 vccd1 vccd1 _12033_/C sky130_fd_sc_hd__nand3_1
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16627__32 vssd1 vssd1 vccd1 vccd1 _16627__32/HI _16693_/A sky130_fd_sc_hd__conb_1
XFILLER_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13982_ _16331_/Q _14039_/B _13989_/C vssd1 vssd1 vccd1 vccd1 _13982_/Y sky130_fd_sc_hd__nand3_1
X_15721_ _15812_/CLK _15721_/D vssd1 vssd1 vccd1 vccd1 _15721_/Q sky130_fd_sc_hd__dfxtp_1
X_12933_ _14060_/A vssd1 vssd1 vccd1 vccd1 _12933_/X sky130_fd_sc_hd__clkbuf_4
X_15652_ _15791_/CLK _15652_/D vssd1 vssd1 vccd1 vccd1 _15652_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _13032_/A _12868_/C vssd1 vssd1 vccd1 vccd1 _12864_/X sky130_fd_sc_hd__or2_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _16423_/Q _14770_/B _14603_/C vssd1 vssd1 vccd1 vccd1 _14612_/B sky130_fd_sc_hd__and3_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _11813_/Y _11814_/X _11810_/C _11811_/C vssd1 vssd1 vccd1 vccd1 _11817_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _16551_/CLK _15583_/D vssd1 vssd1 vccd1 vccd1 _15583_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12793_/Y _12788_/C _12790_/Y _12800_/A vssd1 vssd1 vccd1 vccd1 _12800_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_42_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11746_ _16015_/Q _11969_/B _11757_/C vssd1 vssd1 vccd1 vccd1 _11752_/A sky130_fd_sc_hd__and3_1
X_14534_ _14532_/Y _14527_/C _14529_/Y _14531_/X vssd1 vssd1 vccd1 vccd1 _14535_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11677_ _11903_/A vssd1 vssd1 vccd1 vccd1 _11717_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14465_ _15034_/A vssd1 vssd1 vccd1 vccd1 _14697_/B sky130_fd_sc_hd__buf_2
X_16204_ _16237_/CLK _16204_/D vssd1 vssd1 vccd1 vccd1 _16204_/Q sky130_fd_sc_hd__dfxtp_1
X_10628_ _10652_/C vssd1 vssd1 vccd1 vccd1 _10658_/C sky130_fd_sc_hd__clkbuf_2
X_13416_ _16252_/Q _13586_/B _13416_/C vssd1 vssd1 vccd1 vccd1 _13426_/A sky130_fd_sc_hd__and3_1
X_14396_ _16391_/Q _14433_/C _14339_/X vssd1 vssd1 vccd1 vccd1 _14398_/B sky130_fd_sc_hd__a21oi_1
XFILLER_128_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16135_ _16555_/Q _16135_/D vssd1 vssd1 vccd1 vccd1 _16135_/Q sky130_fd_sc_hd__dfxtp_1
X_13347_ _13354_/A _13347_/B _13347_/C vssd1 vssd1 vccd1 vccd1 _13348_/A sky130_fd_sc_hd__and3_1
X_10559_ _15838_/Q _10652_/B _10559_/C vssd1 vssd1 vccd1 vccd1 _10567_/A sky130_fd_sc_hd__and3_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13278_ _13279_/B _13279_/C _13279_/A vssd1 vssd1 vccd1 vccd1 _13280_/B sky130_fd_sc_hd__a21o_1
X_16066_ _16118_/CLK _16066_/D vssd1 vssd1 vccd1 vccd1 _16066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12229_ _12227_/Y _12222_/C _12224_/Y _12234_/A vssd1 vssd1 vccd1 vccd1 _12234_/B
+ sky130_fd_sc_hd__a211oi_1
X_15017_ _16489_/Q _15055_/C _14906_/X vssd1 vssd1 vccd1 vccd1 _15019_/B sky130_fd_sc_hd__a21oi_1
XFILLER_130_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07770_ _07774_/A vssd1 vssd1 vccd1 vccd1 _07770_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15919_ _15365_/A _15919_/D vssd1 vssd1 vccd1 vccd1 _15919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09440_ _09299_/X _09436_/B _09439_/Y vssd1 vssd1 vccd1 vccd1 _15622_/D sky130_fd_sc_hd__o21a_1
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09371_ _15612_/Q _09416_/B _09371_/C vssd1 vssd1 vccd1 vccd1 _09377_/A sky130_fd_sc_hd__and3_1
XFILLER_80_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08322_ _08143_/A _08143_/B _08321_/Y vssd1 vssd1 vccd1 vccd1 _08345_/A sky130_fd_sc_hd__a21o_1
X_08253_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08275_/A sky130_fd_sc_hd__xnor2_4
XFILLER_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08184_ _12307_/A _07964_/B _07963_/B vssd1 vssd1 vccd1 vccd1 _08186_/C sky130_fd_sc_hd__o21a_1
XFILLER_119_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07968_ _11908_/A _07968_/B vssd1 vssd1 vccd1 vccd1 _08191_/B sky130_fd_sc_hd__xnor2_4
XFILLER_68_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09707_ _10618_/A vssd1 vssd1 vccd1 vccd1 _09707_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07899_ _09987_/C _08296_/B vssd1 vssd1 vccd1 vccd1 _07900_/B sky130_fd_sc_hd__xnor2_2
XFILLER_71_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09638_ _09632_/C _09633_/C _09635_/Y _09642_/A vssd1 vssd1 vccd1 vccd1 _09642_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_71_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09569_ _09524_/X _09567_/B _09568_/Y vssd1 vssd1 vccd1 vccd1 _15648_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11600_ _15995_/Q _11654_/B _11607_/C vssd1 vssd1 vccd1 vccd1 _11600_/X sky130_fd_sc_hd__and3_1
X_12580_ _12580_/A _12580_/B vssd1 vssd1 vccd1 vccd1 _12581_/B sky130_fd_sc_hd__nor2_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11531_ _11525_/C _11526_/C _11528_/Y _11529_/X vssd1 vssd1 vccd1 vccd1 _11532_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14250_ _16371_/Q _14260_/C _14029_/X vssd1 vssd1 vccd1 vccd1 _14250_/Y sky130_fd_sc_hd__a21oi_1
X_11462_ _11520_/A _11462_/B _11467_/A vssd1 vssd1 vccd1 vccd1 _15974_/D sky130_fd_sc_hd__nor3_1
XFILLER_137_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13201_ _13201_/A _13201_/B vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__nor2_1
X_10413_ _10411_/A _10411_/B _10412_/X vssd1 vssd1 vccd1 vccd1 _15810_/D sky130_fd_sc_hd__a21oi_1
XFILLER_139_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14181_ _14175_/C _14176_/C _14178_/Y _14179_/X vssd1 vssd1 vccd1 vccd1 _14182_/C
+ sky130_fd_sc_hd__a211o_1
X_11393_ _11393_/A vssd1 vssd1 vccd1 vccd1 _15965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13132_ _13132_/A vssd1 vssd1 vccd1 vccd1 _16210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10344_ _10337_/C _10338_/C _10341_/Y _10342_/X vssd1 vssd1 vccd1 vccd1 _10345_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_124_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _13058_/Y _13059_/X _13062_/Y _13056_/C vssd1 vssd1 vccd1 vccd1 _13065_/B
+ sky130_fd_sc_hd__o211ai_1
X_10275_ _10220_/X _10268_/B _10271_/B _10274_/Y vssd1 vssd1 vccd1 vccd1 _15784_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12014_ _12183_/A _12018_/C vssd1 vssd1 vccd1 vccd1 _12014_/X sky130_fd_sc_hd__or2_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16753_ _16753_/A _07771_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13965_ _16330_/Q _14185_/B _13966_/C vssd1 vssd1 vccd1 vccd1 _13965_/X sky130_fd_sc_hd__and3_1
XFILLER_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15704_ _15812_/CLK _15704_/D vssd1 vssd1 vccd1 vccd1 _15704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12916_ _16181_/Q _13082_/B _12916_/C vssd1 vssd1 vccd1 vccd1 _12925_/B sky130_fd_sc_hd__and3_1
XFILLER_73_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13896_ _13896_/A _13896_/B _13896_/C vssd1 vssd1 vccd1 vccd1 _13897_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15635_ _15791_/CLK _15635_/D vssd1 vssd1 vccd1 vccd1 _15635_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12847_/A _12847_/B _12847_/C vssd1 vssd1 vccd1 vccd1 _12848_/A sky130_fd_sc_hd__and3_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15566_ _15812_/CLK _15566_/D vssd1 vssd1 vccd1 vccd1 _15566_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _16161_/Q _13009_/B _12778_/C vssd1 vssd1 vccd1 vccd1 _12778_/Y sky130_fd_sc_hd__nand3_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14517_ _14514_/Y _14516_/X _14511_/C _14512_/C vssd1 vssd1 vccd1 vccd1 _14519_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_147_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11729_ _16013_/Q _11950_/B _11729_/C vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__and3_1
X_15497_ _16551_/CLK _15497_/D vssd1 vssd1 vccd1 vccd1 _15497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14448_ _16399_/Q _14486_/C _14339_/X vssd1 vssd1 vccd1 vccd1 _14450_/B sky130_fd_sc_hd__a21oi_1
XFILLER_116_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14379_ _16389_/Q _14380_/C _14265_/X vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__a21oi_1
X_16118_ _16118_/CLK _16118_/D vssd1 vssd1 vccd1 vccd1 _16118_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08940_ _08940_/A _08940_/B _08940_/C vssd1 vssd1 vccd1 vccd1 _08941_/A sky130_fd_sc_hd__and3_1
X_16049_ _16118_/CLK _16049_/D vssd1 vssd1 vccd1 vccd1 _16049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08871_ _08869_/A _08869_/B _08870_/X vssd1 vssd1 vccd1 vccd1 _15502_/D sky130_fd_sc_hd__a21oi_1
XFILLER_97_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ _07824_/A vssd1 vssd1 vccd1 vccd1 _07822_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ _09423_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09423_/X sky130_fd_sc_hd__or2_1
XFILLER_80_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09354_ _09354_/A _09354_/B vssd1 vssd1 vccd1 vccd1 _15605_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08305_ _08314_/A _08314_/B vssd1 vssd1 vccd1 vccd1 _08306_/B sky130_fd_sc_hd__xor2_2
X_09285_ _15262_/B vssd1 vssd1 vccd1 vccd1 _09472_/B sky130_fd_sc_hd__clkbuf_2
X_08236_ _08237_/A _08237_/B vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__or2_4
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08167_ _16607_/Q _08167_/B vssd1 vssd1 vccd1 vccd1 _08167_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08098_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08292_/B sky130_fd_sc_hd__xor2_2
XFILLER_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10060_ _10060_/A vssd1 vssd1 vccd1 vccd1 _10271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10962_ _15905_/Q _10970_/C _10905_/X vssd1 vssd1 vccd1 vccd1 _10962_/Y sky130_fd_sc_hd__a21oi_1
X_13750_ _14308_/A vssd1 vssd1 vccd1 vccd1 _13750_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12701_ _12868_/A _12701_/B _12701_/C vssd1 vssd1 vccd1 vccd1 _12702_/C sky130_fd_sc_hd__or3_1
X_10893_ _15895_/Q _10934_/C _10673_/X vssd1 vssd1 vccd1 vccd1 _10896_/B sky130_fd_sc_hd__a21oi_1
X_13681_ _16290_/Q _13684_/C _13570_/X vssd1 vssd1 vccd1 vccd1 _13681_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15420_ _16221_/Q _16220_/Q _16219_/Q _15416_/X vssd1 vssd1 vccd1 vccd1 _16598_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12632_ _12653_/A _12632_/B _12636_/B vssd1 vssd1 vccd1 vccd1 _16139_/D sky130_fd_sc_hd__nor3_1
X_15351_ _15349_/A _15349_/B _15350_/X vssd1 vssd1 vccd1 vccd1 _16547_/D sky130_fd_sc_hd__a21oi_1
X_12563_ _12559_/Y _12561_/X _12562_/Y _12557_/C vssd1 vssd1 vccd1 vccd1 _12565_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_8_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _11536_/C vssd1 vssd1 vccd1 vccd1 _11551_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14302_ _16378_/Q _14464_/B _14303_/C vssd1 vssd1 vccd1 vccd1 _14302_/X sky130_fd_sc_hd__and3_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15282_ _15282_/A _16702_/A _15282_/C vssd1 vssd1 vccd1 vccd1 _15283_/C sky130_fd_sc_hd__nor3_1
X_12494_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12726_/B sky130_fd_sc_hd__buf_2
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11445_ _11445_/A _11452_/B vssd1 vssd1 vccd1 vccd1 _11447_/A sky130_fd_sc_hd__or2_1
X_14233_ _14256_/A _14233_/B _14233_/C vssd1 vssd1 vccd1 vccd1 _14234_/A sky130_fd_sc_hd__and3_1
XFILLER_125_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14164_ _14164_/A vssd1 vssd1 vccd1 vccd1 _16357_/D sky130_fd_sc_hd__clkbuf_1
X_11376_ _15963_/Q _11495_/B _11381_/C vssd1 vssd1 vccd1 vccd1 _11376_/Y sky130_fd_sc_hd__nand3_1
XFILLER_125_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10327_ _10578_/A vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__buf_2
XFILLER_98_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13115_ _13131_/A _13115_/B _13115_/C vssd1 vssd1 vccd1 vccd1 _13116_/A sky130_fd_sc_hd__and3_1
X_14095_ _14095_/A vssd1 vssd1 vccd1 vccd1 _14318_/B sky130_fd_sc_hd__clkbuf_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _16200_/Q _13053_/C _12879_/X vssd1 vssd1 vccd1 vccd1 _13049_/B sky130_fd_sc_hd__a21o_1
X_10258_ _10338_/A _10258_/B _10258_/C vssd1 vssd1 vccd1 vccd1 _10259_/A sky130_fd_sc_hd__and3_1
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10189_ _15773_/Q _10190_/C _09813_/X vssd1 vssd1 vccd1 vccd1 _10189_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14997_ _14994_/Y _15003_/A _14996_/Y _14992_/C vssd1 vssd1 vccd1 vccd1 _14999_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16736_ _16736_/A _07842_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
XFILLER_81_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13948_ _16327_/Q _13948_/B _13958_/C vssd1 vssd1 vccd1 vccd1 _13953_/A sky130_fd_sc_hd__and3_1
XFILLER_35_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13879_ _13879_/A _13883_/C vssd1 vssd1 vccd1 vccd1 _13879_/X sky130_fd_sc_hd__or2_1
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15618_ _15791_/CLK _15618_/D vssd1 vssd1 vccd1 vccd1 _15618_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16598_ _16607_/CLK _16598_/D vssd1 vssd1 vccd1 vccd1 _16598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15549_ _16551_/CLK _15549_/D vssd1 vssd1 vccd1 vccd1 _15549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09070_ _15551_/Q _09192_/B _09070_/C vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__and3_1
XFILLER_148_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08021_ _10178_/C _08149_/B vssd1 vssd1 vccd1 vccd1 _08022_/B sky130_fd_sc_hd__xnor2_2
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09972_ _10016_/A _09972_/B vssd1 vssd1 vccd1 vccd1 _09973_/B sky130_fd_sc_hd__and2_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08923_ _09125_/A vssd1 vssd1 vccd1 vccd1 _08923_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08854_ _08854_/A vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07805_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07805_/Y sky130_fd_sc_hd__inv_2
X_08785_ _08780_/B _08783_/B _08698_/X vssd1 vssd1 vccd1 vccd1 _08791_/C sky130_fd_sc_hd__o21a_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09406_ _09497_/A _09406_/B _09412_/A vssd1 vssd1 vccd1 vccd1 _15616_/D sky130_fd_sc_hd__nor3_1
XFILLER_53_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09337_ _09336_/X _09335_/Y _10017_/A vssd1 vssd1 vccd1 vccd1 _09337_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09268_ _09265_/Y _09276_/A _09261_/C _09262_/C vssd1 vssd1 vccd1 vccd1 _09270_/B
+ sky130_fd_sc_hd__o211a_1
X_08219_ _08372_/A _08372_/B vssd1 vssd1 vccd1 vccd1 _08220_/B sky130_fd_sc_hd__xor2_4
X_09199_ _10065_/A _09204_/C vssd1 vssd1 vccd1 vccd1 _09199_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _11246_/C vssd1 vssd1 vccd1 vccd1 _11253_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11161_ _15933_/Q _11381_/B _11161_/C vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__and3_1
XFILLER_107_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10112_ _10112_/A vssd1 vssd1 vccd1 vccd1 _10322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11092_ _12225_/A vssd1 vssd1 vccd1 vccd1 _11322_/B sky130_fd_sc_hd__buf_2
XFILLER_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10043_ _15747_/Q _10051_/C _10003_/B vssd1 vssd1 vccd1 vccd1 _10043_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14920_ _14914_/C _14915_/C _14917_/Y _14918_/X vssd1 vssd1 vccd1 vccd1 _14921_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14851_ _14851_/A vssd1 vssd1 vccd1 vccd1 _14851_/X sky130_fd_sc_hd__buf_2
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _13800_/Y _13796_/C _13798_/Y _13799_/X vssd1 vssd1 vccd1 vccd1 _13803_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14782_ _14782_/A vssd1 vssd1 vccd1 vccd1 _16450_/D sky130_fd_sc_hd__clkbuf_1
X_11994_ _16051_/Q _12218_/B _12002_/C vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__and3_1
XFILLER_56_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16521_ _16595_/CLK _16521_/D vssd1 vssd1 vccd1 vccd1 _16521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13733_ _13733_/A _13733_/B _13733_/C vssd1 vssd1 vccd1 vccd1 _13734_/C sky130_fd_sc_hd__nand3_1
X_10945_ _10981_/A _10945_/B _10945_/C vssd1 vssd1 vccd1 vccd1 _10946_/A sky130_fd_sc_hd__and3_1
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ input11/X _16452_/D vssd1 vssd1 vccd1 vccd1 _16452_/Q sky130_fd_sc_hd__dfxtp_2
X_13664_ _16287_/Q _13709_/C _13495_/X vssd1 vssd1 vccd1 vccd1 _13666_/B sky130_fd_sc_hd__a21oi_1
XFILLER_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10876_ input6/X vssd1 vssd1 vccd1 vccd1 _12009_/A sky130_fd_sc_hd__buf_2
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15403_ _15409_/A vssd1 vssd1 vccd1 vccd1 _15403_/X sky130_fd_sc_hd__buf_2
X_12615_ _12612_/Y _12613_/X _12614_/Y _12610_/C vssd1 vssd1 vccd1 vccd1 _12617_/B
+ sky130_fd_sc_hd__o211ai_1
X_16383_ _16389_/CLK _16383_/D vssd1 vssd1 vccd1 vccd1 _16383_/Q sky130_fd_sc_hd__dfxtp_1
X_13595_ _13595_/A _13595_/B vssd1 vssd1 vccd1 vccd1 _13600_/C sky130_fd_sc_hd__nor2_1
X_15334_ _16549_/Q _15335_/C _09364_/B vssd1 vssd1 vccd1 vccd1 _15337_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12546_ _12543_/Y _12545_/X _12540_/C _12541_/C vssd1 vssd1 vccd1 vccd1 _12548_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15265_ _15333_/A _15265_/B _15269_/B vssd1 vssd1 vccd1 vccd1 _16529_/D sky130_fd_sc_hd__nor3_1
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ _16119_/Q _12516_/C _12368_/X vssd1 vssd1 vccd1 vccd1 _12479_/B sky130_fd_sc_hd__a21oi_1
XFILLER_144_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_4 _13886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _14217_/B _14217_/C _14108_/X vssd1 vssd1 vccd1 vccd1 _14218_/B sky130_fd_sc_hd__o21ai_1
X_11428_ _15970_/Q _11488_/B _11436_/C vssd1 vssd1 vccd1 vccd1 _11428_/Y sky130_fd_sc_hd__nand3_1
X_15196_ _15193_/Y _15194_/X _15195_/Y _15191_/C vssd1 vssd1 vccd1 vccd1 _15198_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11359_ _15962_/Q _11359_/B _11361_/C vssd1 vssd1 vccd1 vccd1 _11359_/X sky130_fd_sc_hd__and3_1
X_14147_ _16356_/Q _14154_/C _13979_/X vssd1 vssd1 vccd1 vccd1 _14147_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14078_ _16346_/Q _14185_/B _14079_/C vssd1 vssd1 vccd1 vccd1 _14078_/X sky130_fd_sc_hd__and3_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _13029_/A _13036_/B vssd1 vssd1 vccd1 vccd1 _13031_/A sky130_fd_sc_hd__or2_1
XFILLER_112_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08570_ _08590_/C vssd1 vssd1 vccd1 vccd1 _08619_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16719_ _16719_/A _07823_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
XFILLER_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09122_ _09038_/X _09124_/C _09039_/X vssd1 vssd1 vccd1 vccd1 _09123_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09053_ _15548_/Q _09053_/B _09057_/C vssd1 vssd1 vccd1 vccd1 _09059_/A sky130_fd_sc_hd__and3_1
X_08004_ _08004_/A _08004_/B vssd1 vssd1 vccd1 vccd1 _08020_/A sky130_fd_sc_hd__xor2_4
XFILLER_116_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09955_ _15729_/Q _09998_/B _09955_/C vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__and3_1
XFILLER_106_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08906_ _15515_/Q _08907_/C _08777_/X vssd1 vssd1 vccd1 vccd1 _08908_/A sky130_fd_sc_hd__a21oi_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09884_/X _09886_/B vssd1 vssd1 vccd1 vccd1 _09886_/X sky130_fd_sc_hd__and2b_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08837_ _08706_/X _08835_/A _08833_/X vssd1 vssd1 vccd1 vccd1 _08838_/B sky130_fd_sc_hd__o21ai_1
XFILLER_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08768_ _08768_/A _08768_/B _08768_/C vssd1 vssd1 vccd1 vccd1 _08769_/C sky130_fd_sc_hd__nand3_1
XFILLER_122_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08699_ _08690_/B _08694_/B _08698_/X vssd1 vssd1 vccd1 vccd1 _08705_/C sky130_fd_sc_hd__o21a_1
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10730_ _10731_/B _10731_/C _10731_/A vssd1 vssd1 vccd1 vccd1 _10732_/B sky130_fd_sc_hd__a21o_1
XFILLER_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10661_ _10661_/A _10661_/B vssd1 vssd1 vccd1 vccd1 _10662_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12400_ _12683_/A vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__clkbuf_2
X_13380_ _13401_/C vssd1 vssd1 vccd1 vccd1 _13416_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10592_ _15845_/Q _10593_/C _10492_/X vssd1 vssd1 vccd1 vccd1 _10592_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _16098_/Q _12493_/B _12332_/C vssd1 vssd1 vccd1 vccd1 _12331_/X sky130_fd_sc_hd__and3_1
XFILLER_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15050_ _16493_/Q _15156_/B _15055_/C vssd1 vssd1 vccd1 vccd1 _15050_/Y sky130_fd_sc_hd__nand3_1
X_12262_ _13392_/A vssd1 vssd1 vccd1 vccd1 _12487_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11213_ _11210_/Y _11219_/A _11212_/Y _11208_/C vssd1 vssd1 vccd1 vccd1 _11215_/B
+ sky130_fd_sc_hd__o211a_1
X_14001_ _14017_/C vssd1 vssd1 vccd1 vccd1 _14024_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12193_ _12226_/C vssd1 vssd1 vccd1 vccd1 _12232_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_150_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11144_ _15931_/Q _11367_/B _11152_/C vssd1 vssd1 vccd1 vccd1 _11144_/X sky130_fd_sc_hd__and3_1
XFILLER_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15952_ _15365_/A _15952_/D vssd1 vssd1 vccd1 vccd1 _15952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11075_ _15922_/Q _11078_/C _11023_/X vssd1 vssd1 vccd1 vccd1 _11075_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10026_ _10038_/C vssd1 vssd1 vccd1 vccd1 _10051_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14903_ _14918_/C vssd1 vssd1 vccd1 vccd1 _14925_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15883_ _16553_/Q _15883_/D vssd1 vssd1 vccd1 vccd1 _15883_/Q sky130_fd_sc_hd__dfxtp_1
X_16672__77 vssd1 vssd1 vccd1 vccd1 _16672__77/HI _16748_/A sky130_fd_sc_hd__conb_1
X_14834_ _14834_/A _14834_/B vssd1 vssd1 vccd1 vccd1 _14839_/C sky130_fd_sc_hd__nor2_1
XFILLER_36_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14765_ _16448_/Q _14882_/B _14770_/C vssd1 vssd1 vccd1 vccd1 _14765_/Y sky130_fd_sc_hd__nand3_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11977_ _16049_/Q _11987_/C _11755_/X vssd1 vssd1 vccd1 vccd1 _11977_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16504_ _16607_/CLK _16504_/D vssd1 vssd1 vccd1 vccd1 _16504_/Q sky130_fd_sc_hd__dfxtp_1
X_13716_ _13717_/B _13717_/C _13546_/X vssd1 vssd1 vccd1 vccd1 _13718_/B sky130_fd_sc_hd__o21ai_1
X_10928_ _15900_/Q _11039_/B _10928_/C vssd1 vssd1 vccd1 vccd1 _10936_/A sky130_fd_sc_hd__and3_1
X_14696_ _16438_/Q _14748_/B _14697_/C vssd1 vssd1 vccd1 vccd1 _14696_/X sky130_fd_sc_hd__and3_1
XFILLER_71_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16435_ _16595_/CLK _16435_/D vssd1 vssd1 vccd1 vccd1 _16435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13647_ _13647_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13649_/B sky130_fd_sc_hd__nor2_1
X_10859_ _11993_/A vssd1 vssd1 vccd1 vccd1 _11084_/B sky130_fd_sc_hd__clkbuf_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16389_/CLK _16366_/D vssd1 vssd1 vccd1 vccd1 _16366_/Q sky130_fd_sc_hd__dfxtp_2
X_13578_ _16275_/Q _13586_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13578_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15317_ _15311_/A _15311_/B _15324_/A vssd1 vssd1 vccd1 vccd1 _15317_/Y sky130_fd_sc_hd__a21oi_1
X_12529_ _12683_/A vssd1 vssd1 vccd1 vccd1 _12653_/A sky130_fd_sc_hd__buf_2
XFILLER_145_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16297_ _16533_/Q _16297_/D vssd1 vssd1 vccd1 vccd1 _16297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15248_ _16527_/Q _15248_/B _15248_/C vssd1 vssd1 vccd1 vccd1 _15248_/Y sky130_fd_sc_hd__nand3_1
XFILLER_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _16516_/Q _15232_/B _15188_/C vssd1 vssd1 vccd1 vccd1 _15184_/A sky130_fd_sc_hd__and3_1
XFILLER_98_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09740_ _15686_/Q _09739_/C _09604_/X vssd1 vssd1 vccd1 vccd1 _09741_/B sky130_fd_sc_hd__a21o_1
XFILLER_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
.ends

