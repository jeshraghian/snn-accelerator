* NGSPICE file created from snn.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

.subckt snn clk in1[0] in1[1] in1[2] in1[3] in1[4] in1[5] in1[6] in1[7] io_oeb[0]
+ io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] reset spike_out[0] spike_out[1] state1[0] state1[1] state1[2] state1[3]
+ state1[4] state1[5] state1[6] state1[7] vccd1 vssd1
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09671_ _15408_/Q _09784_/B _09671_/C vssd1 vssd1 vccd1 vccd1 _09671_/X sky130_fd_sc_hd__and3_1
XFILLER_95_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08622_ _15247_/Q _10939_/C _08622_/C vssd1 vssd1 vccd1 vccd1 _08622_/X sky130_fd_sc_hd__and3_1
XFILLER_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08553_ _08611_/A _08553_/B _08557_/A vssd1 vssd1 vccd1 vccd1 _15235_/D sky130_fd_sc_hd__nor3_1
XFILLER_82_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08484_ _12713_/A vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__buf_4
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ _15319_/Q _09334_/B _09105_/C vssd1 vssd1 vccd1 vccd1 _09105_/Y sky130_fd_sc_hd__nand3_1
XFILLER_148_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ _09036_/A _09036_/B _09036_/C vssd1 vssd1 vccd1 vccd1 _09037_/C sky130_fd_sc_hd__nand3_1
XFILLER_89_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09938_ _10114_/A vssd1 vssd1 vccd1 vccd1 _09977_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09869_ _10736_/A vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11900_ _12129_/A vssd1 vssd1 vccd1 vccd1 _11941_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12880_ _12934_/A _12880_/B _12884_/A vssd1 vssd1 vccd1 vccd1 _15909_/D sky130_fd_sc_hd__nor3_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11829_/Y _11824_/C _11836_/A _11828_/Y vssd1 vssd1 vccd1 vccd1 _11836_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14551_/B _14551_/C _14551_/A vssd1 vssd1 vccd1 vccd1 _14552_/B sky130_fd_sc_hd__a21o_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _15733_/Q _11938_/B _11767_/C vssd1 vssd1 vccd1 vccd1 _11762_/Y sky130_fd_sc_hd__nand3_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13507_/A _13499_/Y _13500_/Y _13495_/C vssd1 vssd1 vccd1 vccd1 _13503_/B
+ sky130_fd_sc_hd__o211a_1
X_10713_ _11634_/A vssd1 vssd1 vccd1 vccd1 _10999_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_14_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14481_/A _14481_/B vssd1 vssd1 vccd1 vccd1 _14481_/Y sky130_fd_sc_hd__nor2_1
X_11693_ _11708_/A _11693_/B _11693_/C vssd1 vssd1 vccd1 vccd1 _11694_/A sky130_fd_sc_hd__and3_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16362_/CLK _16220_/D vssd1 vssd1 vccd1 vccd1 _16220_/Q sky130_fd_sc_hd__dfxtp_1
X_13432_ _13430_/X _13431_/Y _13427_/B _13428_/C vssd1 vssd1 vccd1 vccd1 _13434_/B
+ sky130_fd_sc_hd__o211ai_1
X_10644_ _15559_/Q _10817_/B _10654_/C vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__and3_1
XFILLER_9_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _16169_/CLK _16151_/D vssd1 vssd1 vccd1 vccd1 _16151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10575_ _10573_/A _10573_/B _10574_/X vssd1 vssd1 vccd1 vccd1 _15546_/D sky130_fd_sc_hd__a21oi_1
X_13363_ _13362_/X _13360_/C _13206_/X vssd1 vssd1 vccd1 vccd1 _13363_/Y sky130_fd_sc_hd__o21ai_1
X_15102_ _16348_/Q _15171_/B _15107_/C vssd1 vssd1 vccd1 vccd1 _15110_/A sky130_fd_sc_hd__and3_1
X_12314_ _12314_/A _12314_/B _12314_/C vssd1 vssd1 vccd1 vccd1 _12315_/C sky130_fd_sc_hd__nand3_1
X_16082_ _16224_/CLK _16082_/D vssd1 vssd1 vccd1 vccd1 _16082_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13294_ _13300_/A _13292_/Y _13293_/Y _13289_/C vssd1 vssd1 vccd1 vccd1 _13296_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15033_ _15039_/A _15032_/Y _15027_/B _15028_/C vssd1 vssd1 vccd1 vccd1 _15035_/B
+ sky130_fd_sc_hd__o211a_1
X_12245_ _12281_/A _12245_/B _12245_/C vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__and3_1
X_12176_ _12174_/Y _12170_/C _12181_/A _12173_/Y vssd1 vssd1 vccd1 vccd1 _12181_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_123_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11127_ _15635_/Q _11136_/C _10897_/X vssd1 vssd1 vccd1 vccd1 _11127_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11058_ _15624_/Q _11289_/B _11058_/C vssd1 vssd1 vccd1 vccd1 _11058_/X sky130_fd_sc_hd__and3_1
X_15935_ _15935_/CLK _15935_/D vssd1 vssd1 vccd1 vccd1 _15935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10009_ _10064_/A _10009_/B _10013_/A vssd1 vssd1 vccd1 vccd1 _15459_/D sky130_fd_sc_hd__nor3_1
XFILLER_37_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15866_ _07603_/A _15866_/D vssd1 vssd1 vccd1 vccd1 _15866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14817_ _14814_/X _14813_/A _14816_/Y vssd1 vssd1 vccd1 vccd1 _16277_/D sky130_fd_sc_hd__o21a_1
X_15797_ _15195_/Q _15797_/D vssd1 vssd1 vccd1 vccd1 _15797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14748_ _14748_/A _14748_/B _14748_/C vssd1 vssd1 vccd1 vccd1 _14749_/A sky130_fd_sc_hd__and3_1
X_14679_ _14679_/A _14679_/B vssd1 vssd1 vccd1 vccd1 _14682_/A sky130_fd_sc_hd__or2_1
XFILLER_20_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ _16358_/CLK _16349_/D vssd1 vssd1 vccd1 vccd1 _16349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07984_ _07984_/A _08177_/A vssd1 vssd1 vccd1 vccd1 _07985_/B sky130_fd_sc_hd__xnor2_2
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09723_ _09724_/B _09724_/C _09724_/A vssd1 vssd1 vccd1 vccd1 _09725_/B sky130_fd_sc_hd__a21o_1
XFILLER_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09654_ _09690_/A _09654_/B _09654_/C vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__and3_1
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08605_ _15260_/Q _15259_/Q _15258_/Q _08604_/X vssd1 vssd1 vccd1 vccd1 _15243_/D
+ sky130_fd_sc_hd__o31a_1
X_09585_ _15394_/Q _09644_/B _09585_/C vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__and3_1
XFILLER_63_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08536_ _08536_/A _08536_/B vssd1 vssd1 vccd1 vccd1 _08540_/C sky130_fd_sc_hd__nor2_1
XFILLER_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08467_ _08467_/A vssd1 vssd1 vccd1 vccd1 _15221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08398_ _08372_/A _08378_/A _08411_/A _08397_/Y vssd1 vssd1 vccd1 vccd1 _08400_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10360_ _10360_/A _10360_/B _10360_/C vssd1 vssd1 vccd1 vccd1 _10361_/C sky130_fd_sc_hd__nand3_1
X_09019_ _14372_/A vssd1 vssd1 vccd1 vccd1 _09019_/X sky130_fd_sc_hd__clkbuf_2
X_10291_ _10312_/C vssd1 vssd1 vccd1 vccd1 _10325_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12030_ _12030_/A _12030_/B _12030_/C vssd1 vssd1 vccd1 vccd1 _12031_/C sky130_fd_sc_hd__nand3_1
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13981_ _16103_/Q _13981_/B _13990_/C vssd1 vssd1 vccd1 vccd1 _13985_/B sky130_fd_sc_hd__nand3_1
XFILLER_120_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15720_ _15794_/CLK _15720_/D vssd1 vssd1 vccd1 vccd1 _15720_/Q sky130_fd_sc_hd__dfxtp_2
X_12932_ _15919_/Q _12968_/C _12767_/X vssd1 vssd1 vccd1 vccd1 _12934_/B sky130_fd_sc_hd__a21oi_1
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15651_ _15655_/CLK _15651_/D vssd1 vssd1 vccd1 vccd1 _15651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12863_ _12869_/B _12863_/B vssd1 vssd1 vccd1 vccd1 _12865_/A sky130_fd_sc_hd__or2_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14601_/X _14600_/Y _14648_/A vssd1 vssd1 vccd1 vccd1 _14602_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _15741_/Q _11986_/B _11814_/C vssd1 vssd1 vccd1 vccd1 _11814_/Y sky130_fd_sc_hd__nand3_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15194_/Q _15582_/D vssd1 vssd1 vccd1 vccd1 _15582_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12791_/X _12792_/Y _12793_/Y _12789_/C vssd1 vssd1 vccd1 vccd1 _12796_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14533_/A _14533_/B vssd1 vssd1 vccd1 vccd1 _14533_/Y sky130_fd_sc_hd__nor2_1
X_11745_ _15732_/Q _11863_/B _11745_/C vssd1 vssd1 vccd1 vccd1 _11745_/X sky130_fd_sc_hd__and3_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464_ _14474_/C vssd1 vssd1 vccd1 vccd1 _14486_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11676_ _11676_/A vssd1 vssd1 vccd1 vccd1 _11689_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16203_ _16204_/CLK _16203_/D vssd1 vssd1 vccd1 vccd1 _16203_/Q sky130_fd_sc_hd__dfxtp_1
X_13415_ _16016_/Q _16015_/Q _16014_/Q _13209_/X vssd1 vssd1 vccd1 vccd1 _15999_/D
+ sky130_fd_sc_hd__o31a_1
X_10627_ _10627_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10628_/B sky130_fd_sc_hd__nor2_1
X_14395_ _14395_/A vssd1 vssd1 vccd1 vccd1 _14395_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16134_ _16143_/CLK _16134_/D vssd1 vssd1 vccd1 vccd1 _16134_/Q sky130_fd_sc_hd__dfxtp_1
X_13346_ _13352_/A _13343_/Y _13345_/Y _13339_/C vssd1 vssd1 vccd1 vccd1 _13348_/B
+ sky130_fd_sc_hd__o211a_1
X_10558_ _10556_/Y _10552_/C _10554_/X _10555_/Y vssd1 vssd1 vccd1 vccd1 _10559_/C
+ sky130_fd_sc_hd__a211o_1
X_16065_ _16075_/CLK _16065_/D vssd1 vssd1 vccd1 vccd1 _16065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13277_ _14080_/B vssd1 vssd1 vccd1 vccd1 _13277_/X sky130_fd_sc_hd__clkbuf_4
X_10489_ _10489_/A vssd1 vssd1 vccd1 vccd1 _15533_/D sky130_fd_sc_hd__clkbuf_1
X_15016_ _15013_/X _15012_/A _15015_/Y vssd1 vssd1 vccd1 vccd1 _16322_/D sky130_fd_sc_hd__o21a_1
X_12228_ _15807_/Q _12228_/B _12228_/C vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__and3_1
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12159_ _15795_/Q _12270_/B _12159_/C vssd1 vssd1 vccd1 vccd1 _12159_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15918_ _15196_/Q _15918_/D vssd1 vssd1 vccd1 vccd1 _15918_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15849_ _15907_/CLK _15849_/D vssd1 vssd1 vccd1 vccd1 _15849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09370_ _09403_/C vssd1 vssd1 vccd1 vccd1 _09411_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_52_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08321_ _08321_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08324_/A sky130_fd_sc_hd__xnor2_2
XFILLER_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08252_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08252_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08183_ _08042_/A _08042_/B _08182_/X vssd1 vssd1 vccd1 vccd1 _08199_/A sky130_fd_sc_hd__a21bo_1
XFILLER_119_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07967_ _16215_/Q _07967_/B vssd1 vssd1 vccd1 vccd1 _07967_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09706_ _09704_/A _09704_/B _09705_/X vssd1 vssd1 vccd1 vccd1 _15411_/D sky130_fd_sc_hd__a21oi_1
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07898_ _15476_/Q vssd1 vssd1 vccd1 vccd1 _10121_/A sky130_fd_sc_hd__inv_2
X_09637_ _09924_/A vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ _09575_/A _09568_/B _09568_/C vssd1 vssd1 vccd1 vccd1 _09569_/A sky130_fd_sc_hd__and3_1
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08519_ _08519_/A _08519_/B _08519_/C vssd1 vssd1 vccd1 vccd1 _08520_/A sky130_fd_sc_hd__and3_1
XFILLER_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ _09496_/X _09498_/Y _09493_/B _09494_/C vssd1 vssd1 vccd1 vccd1 _09501_/B
+ sky130_fd_sc_hd__o211ai_1
X_11530_ _11528_/Y _11523_/C _11525_/X _11527_/Y vssd1 vssd1 vccd1 vccd1 _11531_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11461_ _11477_/A _11461_/B _11461_/C vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__and3_1
XFILLER_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13200_ _13198_/A _13198_/B _13199_/X vssd1 vssd1 vccd1 vccd1 _15960_/D sky130_fd_sc_hd__a21oi_1
X_10412_ _10426_/C vssd1 vssd1 vccd1 vccd1 _10434_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11392_ _15676_/Q _11431_/C _11336_/X vssd1 vssd1 vccd1 vccd1 _11394_/B sky130_fd_sc_hd__a21oi_1
X_14180_ _14180_/A _14180_/B vssd1 vssd1 vccd1 vccd1 _14180_/X sky130_fd_sc_hd__or2_1
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _14261_/A vssd1 vssd1 vccd1 vccd1 _14395_/A sky130_fd_sc_hd__buf_4
X_10343_ _10342_/B _10342_/C _10172_/X vssd1 vssd1 vccd1 vccd1 _10344_/C sky130_fd_sc_hd__o21ai_1
XFILLER_109_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10274_ _10353_/A _10274_/B _10279_/B vssd1 vssd1 vccd1 vccd1 _15500_/D sky130_fd_sc_hd__nor3_1
X_13062_ _13069_/A _13062_/B _13062_/C vssd1 vssd1 vccd1 vccd1 _13063_/A sky130_fd_sc_hd__and3_1
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12013_ _12011_/A _12011_/B _12012_/X vssd1 vssd1 vccd1 vccd1 _15771_/D sky130_fd_sc_hd__a21oi_1
XFILLER_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_2_0_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_7_clk/A sky130_fd_sc_hd__clkbuf_16
XFILLER_47_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13964_ _14054_/A _13964_/B vssd1 vssd1 vccd1 vccd1 _13964_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _15794_/CLK _15703_/D vssd1 vssd1 vccd1 vccd1 _15703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12915_ _15916_/Q _12914_/C _10970_/C vssd1 vssd1 vccd1 vccd1 _12916_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13895_ _13895_/A _13895_/B vssd1 vssd1 vccd1 vccd1 _13895_/Y sky130_fd_sc_hd__nor2_1
X_15634_ _15194_/Q _15634_/D vssd1 vssd1 vccd1 vccd1 _15634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12846_ _15905_/Q _12854_/C _12616_/X vssd1 vssd1 vccd1 vccd1 _12846_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _15655_/CLK _15565_/D vssd1 vssd1 vccd1 vccd1 _15565_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12996_/B sky130_fd_sc_hd__buf_2
XFILLER_42_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14510_/B _14511_/C _14520_/A _14514_/Y vssd1 vssd1 vccd1 vccd1 _14520_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _11727_/B _11727_/C _11615_/X vssd1 vssd1 vccd1 vccd1 _11729_/C sky130_fd_sc_hd__o21ai_1
X_15496_ _15224_/Q _15496_/D vssd1 vssd1 vccd1 vccd1 _15496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14447_ _16196_/Q _14566_/B _14447_/C vssd1 vssd1 vccd1 vccd1 _14447_/X sky130_fd_sc_hd__and3_1
X_11659_ _11665_/A _11656_/Y _11658_/Y _11653_/C vssd1 vssd1 vccd1 vccd1 _11661_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14378_ _16183_/Q _14403_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14381_/B sky130_fd_sc_hd__a21oi_1
XFILLER_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16117_ _16119_/CLK _16117_/D vssd1 vssd1 vccd1 vccd1 _16117_/Q sky130_fd_sc_hd__dfxtp_2
X_13329_ _13327_/X _13328_/Y _13324_/B _13325_/C vssd1 vssd1 vccd1 vccd1 _13331_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 _15584_/CLK sky130_fd_sc_hd__clkbuf_2
X_16048_ _16060_/CLK _16048_/D vssd1 vssd1 vccd1 vccd1 _16048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08870_ _08878_/A _08870_/B _08870_/C vssd1 vssd1 vccd1 vccd1 _08871_/A sky130_fd_sc_hd__and3_1
XFILLER_123_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07821_ _07821_/A _07821_/B vssd1 vssd1 vccd1 vccd1 _07822_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07752_ _07752_/A _07752_/B vssd1 vssd1 vccd1 vccd1 _07754_/B sky130_fd_sc_hd__xor2_4
XFILLER_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07683_ _14099_/B vssd1 vssd1 vccd1 vccd1 _14364_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09422_ _09422_/A vssd1 vssd1 vccd1 vccd1 _15367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09353_ _09353_/A _09353_/B _09357_/B vssd1 vssd1 vccd1 vccd1 _15357_/D sky130_fd_sc_hd__nor3_1
XFILLER_80_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08304_ _08304_/A _08352_/A vssd1 vssd1 vccd1 vccd1 _08343_/A sky130_fd_sc_hd__xnor2_2
X_09284_ _15348_/Q _09290_/C _09166_/X vssd1 vssd1 vccd1 vccd1 _09284_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ _08103_/A _08103_/B _08234_/Y vssd1 vssd1 vccd1 vccd1 _08239_/A sky130_fd_sc_hd__a21o_1
X_08166_ _08429_/C _08166_/B vssd1 vssd1 vccd1 vccd1 _08166_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08097_ _08238_/A _08097_/B vssd1 vssd1 vccd1 vccd1 _08234_/A sky130_fd_sc_hd__nand2_2
XFILLER_107_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08999_ _08999_/A _08999_/B _08999_/C vssd1 vssd1 vccd1 vccd1 _09000_/A sky130_fd_sc_hd__and3_1
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10961_ _10961_/A vssd1 vssd1 vccd1 vccd1 _15607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12700_ _12699_/B _12699_/C _12472_/X vssd1 vssd1 vccd1 vccd1 _12701_/C sky130_fd_sc_hd__o21ai_1
X_13680_ _16048_/Q _14074_/B _13686_/C vssd1 vssd1 vccd1 vccd1 _13683_/B sky130_fd_sc_hd__nand3_1
X_10892_ _10890_/Y _10886_/C _10888_/X _10889_/Y vssd1 vssd1 vccd1 vccd1 _10893_/C
+ sky130_fd_sc_hd__a211o_1
X_12631_ _12631_/A vssd1 vssd1 vccd1 vccd1 _12631_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15350_ _15356_/CLK _15350_/D vssd1 vssd1 vccd1 vccd1 _15350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ _15859_/Q _12793_/B _12568_/C vssd1 vssd1 vccd1 vccd1 _12562_/Y sky130_fd_sc_hd__nand3_1
X_14301_ _16167_/Q _14299_/C _14300_/X vssd1 vssd1 vccd1 vccd1 _14301_/Y sky130_fd_sc_hd__a21oi_1
X_11513_ _15695_/Q _11518_/C _11512_/X vssd1 vssd1 vccd1 vccd1 _11515_/C sky130_fd_sc_hd__a21o_1
X_15281_ _15282_/CLK _15281_/D vssd1 vssd1 vccd1 vccd1 _15281_/Q sky130_fd_sc_hd__dfxtp_1
X_12493_ _15849_/Q _12500_/C _12377_/X vssd1 vssd1 vccd1 vccd1 _12493_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14232_ _14227_/Y _14230_/X _14231_/Y vssd1 vssd1 vccd1 vccd1 _16148_/D sky130_fd_sc_hd__o21a_1
X_11444_ _15683_/Q vssd1 vssd1 vccd1 vccd1 _11457_/C sky130_fd_sc_hd__inv_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14163_ _14163_/A vssd1 vssd1 vccd1 vccd1 _14979_/A sky130_fd_sc_hd__buf_4
X_11375_ _15673_/Q _11374_/C _11199_/X vssd1 vssd1 vccd1 vccd1 _11376_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13114_ _13149_/A _13114_/B _13114_/C vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__and3_1
X_10326_ _15510_/Q _10331_/C _10269_/X vssd1 vssd1 vccd1 vccd1 _10326_/Y sky130_fd_sc_hd__a21oi_1
X_14094_ _16123_/Q _14099_/C _14270_/A vssd1 vssd1 vccd1 vccd1 _14094_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _15939_/Q _13045_/B _13051_/C vssd1 vssd1 vccd1 vccd1 _13048_/B sky130_fd_sc_hd__nand3_1
X_10257_ _10253_/X _10254_/Y _10256_/Y _10251_/C vssd1 vssd1 vccd1 vccd1 _10259_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ _10188_/A _10188_/B _10188_/C vssd1 vssd1 vccd1 vccd1 _10189_/C sky130_fd_sc_hd__nand3_1
XFILLER_66_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14996_ _14996_/A _14996_/B vssd1 vssd1 vccd1 vccd1 _14998_/A sky130_fd_sc_hd__or2_1
XFILLER_19_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13947_ _13952_/A _13946_/Y _13942_/B _13943_/C vssd1 vssd1 vccd1 vccd1 _13949_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13878_ _14291_/A vssd1 vssd1 vccd1 vccd1 _14587_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15617_ _15194_/Q _15617_/D vssd1 vssd1 vccd1 vccd1 _15617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12829_ _12829_/A _12829_/B _12829_/C vssd1 vssd1 vccd1 vccd1 _12830_/C sky130_fd_sc_hd__nand3_1
X_15548_ _15656_/CLK _15548_/D vssd1 vssd1 vccd1 vccd1 _15548_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15479_ _15483_/CLK _15479_/D vssd1 vssd1 vccd1 vccd1 _15479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _08020_/A _08020_/B vssd1 vssd1 vccd1 vccd1 _08021_/B sky130_fd_sc_hd__nor2_2
XFILLER_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ _09971_/A vssd1 vssd1 vccd1 vccd1 _15453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08922_ _08919_/X _08921_/Y _08916_/B _08917_/C vssd1 vssd1 vccd1 vccd1 _08924_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_130_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08853_ _15282_/Q _08853_/B _08859_/C vssd1 vssd1 vccd1 vccd1 _08856_/B sky130_fd_sc_hd__nand3_1
XFILLER_111_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07804_ _15845_/Q _08049_/B vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__xnor2_2
XFILLER_57_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08784_ _08783_/B _08783_/C _08726_/X vssd1 vssd1 vccd1 vccd1 _08785_/C sky130_fd_sc_hd__o21ai_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07735_ _08109_/A _07735_/B vssd1 vssd1 vccd1 vccd1 _07738_/B sky130_fd_sc_hd__xnor2_1
XFILLER_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07666_ _07666_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09405_ _15366_/Q _09411_/C _09404_/X vssd1 vssd1 vccd1 vccd1 _09405_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07597_ input9/X vssd1 vssd1 vccd1 vccd1 _13930_/A sky130_fd_sc_hd__buf_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09336_ _09334_/Y _09330_/C _09332_/X _09333_/Y vssd1 vssd1 vccd1 vccd1 _09337_/C
+ sky130_fd_sc_hd__a211o_1
X_09267_ _09288_/A _09267_/B _09267_/C vssd1 vssd1 vccd1 vccd1 _09268_/A sky130_fd_sc_hd__and3_1
XFILLER_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _08218_/A _08218_/B vssd1 vssd1 vccd1 vccd1 _08219_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09198_ _09222_/C vssd1 vssd1 vccd1 vccd1 _09236_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08149_ _07893_/A _07893_/B _08148_/Y vssd1 vssd1 vccd1 vccd1 _08264_/B sky130_fd_sc_hd__o21a_1
XFILLER_134_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11160_ _15640_/Q _11198_/C _11047_/X vssd1 vssd1 vccd1 vccd1 _11162_/B sky130_fd_sc_hd__a21oi_1
XFILLER_122_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ _10111_/A _10111_/B vssd1 vssd1 vccd1 vccd1 _10115_/C sky130_fd_sc_hd__nor2_1
X_11091_ _11204_/A _11094_/C vssd1 vssd1 vccd1 vccd1 _11091_/X sky130_fd_sc_hd__or2_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10042_ _10064_/A _10042_/B _10047_/B vssd1 vssd1 vccd1 vccd1 _15464_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14850_ _14766_/X _14853_/C _14808_/X vssd1 vssd1 vccd1 vccd1 _14851_/B sky130_fd_sc_hd__o21ai_1
XFILLER_29_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13801_ _16068_/Q _13801_/B _13805_/C vssd1 vssd1 vccd1 vccd1 _13801_/Y sky130_fd_sc_hd__nand3_1
X_14781_ _14980_/A vssd1 vssd1 vccd1 vccd1 _14941_/B sky130_fd_sc_hd__clkbuf_2
X_11993_ _12277_/A vssd1 vssd1 vccd1 vccd1 _12223_/B sky130_fd_sc_hd__clkbuf_2
X_13732_ _16057_/Q _13738_/C _13526_/X vssd1 vssd1 vccd1 vccd1 _13734_/C sky130_fd_sc_hd__a21o_1
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10944_ _10960_/A _10944_/B _10944_/C vssd1 vssd1 vccd1 vccd1 _10945_/A sky130_fd_sc_hd__and3_1
XFILLER_45_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13663_ _13662_/B _13662_/C _13562_/X vssd1 vssd1 vccd1 vccd1 _13664_/C sky130_fd_sc_hd__o21ai_1
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10875_ _10931_/A _10875_/B _10879_/A vssd1 vssd1 vccd1 vccd1 _15594_/D sky130_fd_sc_hd__nor3_1
XFILLER_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15402_ _15484_/CLK _15402_/D vssd1 vssd1 vccd1 vccd1 _15402_/Q sky130_fd_sc_hd__dfxtp_1
X_12614_ _12614_/A vssd1 vssd1 vccd1 vccd1 _15867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13594_ _13592_/Y _13587_/C _13589_/X _13590_/Y vssd1 vssd1 vccd1 vccd1 _13595_/C
+ sky130_fd_sc_hd__a211o_1
X_15333_ _15333_/CLK _15333_/D vssd1 vssd1 vccd1 vccd1 _15333_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12545_ _12545_/A vssd1 vssd1 vccd1 vccd1 _15856_/D sky130_fd_sc_hd__clkbuf_1
X_15264_ _15274_/CLK _15264_/D vssd1 vssd1 vccd1 vccd1 _15264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12476_ _15853_/Q _15852_/Q _15851_/Q _12418_/X vssd1 vssd1 vccd1 vccd1 _15845_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_144_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14215_ _14434_/A vssd1 vssd1 vccd1 vccd1 _14304_/A sky130_fd_sc_hd__clkbuf_2
X_11427_ _15680_/Q _11601_/B _11431_/C vssd1 vssd1 vccd1 vccd1 _11427_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_5 state1[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15195_ _15194_/Q _15195_/D vssd1 vssd1 vccd1 vccd1 _15195_/Q sky130_fd_sc_hd__dfxtp_4
X_14146_ _14321_/A _14146_/B vssd1 vssd1 vccd1 vccd1 _14146_/Y sky130_fd_sc_hd__nor2_1
X_11358_ _11365_/A _11358_/B _11358_/C vssd1 vssd1 vccd1 vccd1 _11359_/A sky130_fd_sc_hd__and3_1
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _10309_/A vssd1 vssd1 vccd1 vccd1 _15506_/D sky130_fd_sc_hd__clkbuf_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14077_ _14077_/A _14077_/B _14077_/C vssd1 vssd1 vccd1 vccd1 _14078_/C sky130_fd_sc_hd__nand3_1
X_11289_ _15660_/Q _11289_/B _11289_/C vssd1 vssd1 vccd1 vccd1 _11289_/X sky130_fd_sc_hd__and3_1
XFILLER_79_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _13026_/A _13026_/B _13027_/X vssd1 vssd1 vccd1 vccd1 _15933_/D sky130_fd_sc_hd__a21oi_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14979_ _14979_/A vssd1 vssd1 vccd1 vccd1 _15135_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09121_ _09128_/A _09119_/Y _09120_/Y _09115_/C vssd1 vssd1 vccd1 vccd1 _09123_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09052_ _15312_/Q _09165_/B _09061_/C vssd1 vssd1 vccd1 vccd1 _09052_/X sky130_fd_sc_hd__and3_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08003_ _13777_/C _07880_/B _07879_/A vssd1 vssd1 vccd1 vccd1 _08205_/A sky130_fd_sc_hd__o21a_2
XFILLER_143_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _09955_/B _09955_/C _09955_/A vssd1 vssd1 vccd1 vccd1 _09956_/B sky130_fd_sc_hd__a21o_1
XFILLER_89_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08905_ _08931_/C vssd1 vssd1 vccd1 vccd1 _08945_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _09883_/B _09883_/C _09884_/X vssd1 vssd1 vccd1 vccd1 _09886_/C sky130_fd_sc_hd__o21ai_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08836_ _08893_/A _08839_/C vssd1 vssd1 vccd1 vccd1 _08836_/X sky130_fd_sc_hd__or2_1
XFILLER_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08767_ input6/X vssd1 vssd1 vccd1 vccd1 _09924_/A sky130_fd_sc_hd__buf_4
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07718_ _15252_/Q vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__clkinv_2
X_08698_ _08698_/A vssd1 vssd1 vccd1 vccd1 _15256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07649_ _15171_/B vssd1 vssd1 vccd1 vccd1 _07649_/X sky130_fd_sc_hd__buf_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ _10660_/A vssd1 vssd1 vccd1 vccd1 _15560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09319_ _09353_/A _09319_/B _09323_/A vssd1 vssd1 vccd1 vccd1 _15352_/D sky130_fd_sc_hd__nor3_1
X_10591_ _15551_/Q _10596_/C _10357_/X vssd1 vssd1 vccd1 vccd1 _10593_/C sky130_fd_sc_hd__a21o_1
X_12330_ _12330_/A vssd1 vssd1 vccd1 vccd1 _15822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12261_ _12261_/A vssd1 vssd1 vccd1 vccd1 _15811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14000_ _13999_/X _13998_/Y _14612_/A vssd1 vssd1 vccd1 vccd1 _14000_/Y sky130_fd_sc_hd__a21oi_1
X_11212_ _15655_/Q _15654_/Q _15653_/Q _10983_/X vssd1 vssd1 vccd1 vccd1 _15647_/D
+ sky130_fd_sc_hd__o31a_1
X_12192_ _15808_/Q _15807_/Q _15806_/Q _12134_/X vssd1 vssd1 vccd1 vccd1 _15800_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_134_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11143_ _15637_/Q _11143_/B _11143_/C vssd1 vssd1 vccd1 vccd1 _11151_/B sky130_fd_sc_hd__and3_1
XFILLER_96_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11074_ _11071_/X _11072_/Y _11073_/Y _11069_/C vssd1 vssd1 vccd1 vccd1 _11076_/B
+ sky130_fd_sc_hd__o211ai_1
X_15951_ _16100_/CLK _15951_/D vssd1 vssd1 vccd1 vccd1 _15951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10025_ _10022_/X _10023_/Y _10024_/Y _10020_/C vssd1 vssd1 vccd1 vccd1 _10027_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_49_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14902_ _16301_/Q _14916_/C _14901_/X vssd1 vssd1 vccd1 vccd1 _14904_/B sky130_fd_sc_hd__a21oi_1
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15882_ _07603_/A _15882_/D vssd1 vssd1 vccd1 vccd1 _15882_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14833_ _16285_/Q _14833_/B _14838_/C vssd1 vssd1 vccd1 vccd1 _14841_/A sky130_fd_sc_hd__and3_1
XFILLER_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14764_ _07675_/X _14757_/A _14760_/B _14763_/Y vssd1 vssd1 vccd1 vccd1 _16265_/D
+ sky130_fd_sc_hd__o31a_1
X_11976_ _11997_/A _11976_/B _11976_/C vssd1 vssd1 vccd1 vccd1 _11977_/A sky130_fd_sc_hd__and3_1
XFILLER_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13715_ _13715_/A vssd1 vssd1 vccd1 vccd1 _14106_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10927_ _10950_/B vssd1 vssd1 vccd1 vccd1 _10963_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14695_ _15169_/A vssd1 vssd1 vccd1 vccd1 _14695_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13646_ _13664_/A _13646_/B _13646_/C vssd1 vssd1 vccd1 vccd1 _13647_/A sky130_fd_sc_hd__and3_1
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10858_ _10858_/A _10858_/B vssd1 vssd1 vccd1 vccd1 _10859_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _16367_/CLK _16365_/D vssd1 vssd1 vccd1 vccd1 _16365_/Q sky130_fd_sc_hd__dfxtp_1
X_13577_ _16030_/Q _13628_/B _13583_/C vssd1 vssd1 vccd1 vccd1 _13580_/B sky130_fd_sc_hd__nand3_1
X_10789_ _10789_/A _10789_/B _10789_/C vssd1 vssd1 vccd1 vccd1 _10790_/A sky130_fd_sc_hd__and3_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15316_ _16317_/CLK _15316_/D vssd1 vssd1 vccd1 vccd1 _15316_/Q sky130_fd_sc_hd__dfxtp_2
X_12528_ _12527_/B _12527_/C _12472_/X vssd1 vssd1 vccd1 vccd1 _12529_/C sky130_fd_sc_hd__o21ai_1
X_16296_ _16317_/CLK _16296_/D vssd1 vssd1 vccd1 vccd1 _16296_/Q sky130_fd_sc_hd__dfxtp_1
X_15247_ _15351_/CLK _15247_/D vssd1 vssd1 vccd1 vccd1 _15247_/Q sky130_fd_sc_hd__dfxtp_1
X_12459_ _12465_/A _12457_/Y _12458_/Y _12454_/C vssd1 vssd1 vccd1 vccd1 _12461_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15178_ _15178_/A _15178_/B vssd1 vssd1 vccd1 vccd1 _15180_/A sky130_fd_sc_hd__or2_1
XFILLER_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14129_ _14208_/A _14129_/B _14132_/B vssd1 vssd1 vccd1 vccd1 _16128_/D sky130_fd_sc_hd__nor3_1
XFILLER_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ _09670_/A vssd1 vssd1 vccd1 vccd1 _15406_/D sky130_fd_sc_hd__clkbuf_1
X_08621_ _08621_/A vssd1 vssd1 vccd1 vccd1 _15245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08552_ _15236_/Q _08794_/B _08560_/C vssd1 vssd1 vccd1 vccd1 _08557_/A sky130_fd_sc_hd__and3_1
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08483_ input2/X vssd1 vssd1 vccd1 vccd1 _12713_/A sky130_fd_sc_hd__buf_2
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09104_ _13534_/A vssd1 vssd1 vccd1 vccd1 _09334_/B sky130_fd_sc_hd__clkbuf_4
X_09035_ _09036_/B _09036_/C _09036_/A vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__a21o_1
XFILLER_117_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09937_ _09935_/A _09935_/B _09936_/X vssd1 vssd1 vccd1 vccd1 _15447_/D sky130_fd_sc_hd__a21oi_1
XFILLER_131_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09868_ _15438_/Q _09874_/C _09693_/X vssd1 vssd1 vccd1 vccd1 _09868_/Y sky130_fd_sc_hd__a21oi_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08819_ _08816_/X _08817_/Y _08818_/Y _08814_/C vssd1 vssd1 vccd1 vccd1 _08821_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_133_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09799_ _09807_/A _09799_/B _09799_/C vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__and3_1
XFILLER_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _11836_/A _11828_/Y _11829_/Y _11824_/C vssd1 vssd1 vccd1 vccd1 _11832_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _15734_/Q _11767_/C _11760_/X vssd1 vssd1 vccd1 vccd1 _11761_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _16014_/Q _13550_/B _13504_/C vssd1 vssd1 vccd1 vccd1 _13500_/Y sky130_fd_sc_hd__nand3_1
X_10712_ _10712_/A vssd1 vssd1 vccd1 vccd1 _15568_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _16204_/Q _14486_/C _14395_/X vssd1 vssd1 vccd1 vccd1 _14482_/B sky130_fd_sc_hd__a21oi_1
X_11692_ _11686_/B _11687_/C _11689_/X _11690_/Y vssd1 vssd1 vccd1 vccd1 _11693_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _16004_/Q _13430_/C _13277_/X vssd1 vssd1 vccd1 vccd1 _13431_/Y sky130_fd_sc_hd__a21oi_1
X_10643_ _15559_/Q _10685_/C _10474_/X vssd1 vssd1 vccd1 vccd1 _10645_/B sky130_fd_sc_hd__a21oi_1
XFILLER_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16150_ _16169_/CLK _16150_/D vssd1 vssd1 vccd1 vccd1 _16150_/Q sky130_fd_sc_hd__dfxtp_1
X_13362_ _13617_/A vssd1 vssd1 vccd1 vccd1 _13362_/X sky130_fd_sc_hd__clkbuf_2
X_10574_ _10629_/A _10577_/C vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__or2_1
X_15101_ _15101_/A vssd1 vssd1 vccd1 vccd1 _16343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12313_ _12314_/B _12314_/C _12314_/A vssd1 vssd1 vccd1 vccd1 _12315_/B sky130_fd_sc_hd__a21o_1
X_16081_ _16224_/CLK _16081_/D vssd1 vssd1 vccd1 vccd1 _16081_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13293_ _15978_/Q _13293_/B _13297_/C vssd1 vssd1 vccd1 vccd1 _13293_/Y sky130_fd_sc_hd__nand3_1
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15032_ _16330_/Q _15036_/C _14988_/X vssd1 vssd1 vccd1 vccd1 _15032_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12244_ _12243_/B _12243_/C _12188_/X vssd1 vssd1 vccd1 vccd1 _12245_/C sky130_fd_sc_hd__o21ai_1
XFILLER_122_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ _12181_/A _12173_/Y _12174_/Y _12170_/C vssd1 vssd1 vccd1 vccd1 _12177_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11126_ _15635_/Q _11244_/B _11136_/C vssd1 vssd1 vccd1 vccd1 _11126_/X sky130_fd_sc_hd__and3_1
XFILLER_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11057_ _11634_/A vssd1 vssd1 vccd1 vccd1 _11289_/B sky130_fd_sc_hd__clkbuf_2
X_15934_ _15196_/Q _15934_/D vssd1 vssd1 vccd1 vccd1 _15934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10008_ _15460_/Q _10239_/B _10016_/C vssd1 vssd1 vccd1 vccd1 _10013_/A sky130_fd_sc_hd__and3_1
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15865_ _07603_/A _15865_/D vssd1 vssd1 vccd1 vccd1 _15865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14816_ _14772_/X _14813_/A _14815_/X vssd1 vssd1 vccd1 vccd1 _14816_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15796_ _15195_/Q _15796_/D vssd1 vssd1 vccd1 vccd1 _15796_/Q sky130_fd_sc_hd__dfxtp_1
X_11959_ _11958_/B _11958_/C _11902_/X vssd1 vssd1 vccd1 vccd1 _11960_/C sky130_fd_sc_hd__o21ai_1
X_14747_ _14747_/A _14747_/B _14747_/C vssd1 vssd1 vccd1 vccd1 _14748_/C sky130_fd_sc_hd__nand3_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14678_ _16250_/Q _14677_/C _14095_/B vssd1 vssd1 vccd1 vccd1 _14679_/B sky130_fd_sc_hd__a21oi_1
X_13629_ _16039_/Q _13634_/C _13526_/X vssd1 vssd1 vccd1 vccd1 _13631_/C sky130_fd_sc_hd__a21o_1
XFILLER_20_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348_ _16364_/CLK _16348_/D vssd1 vssd1 vccd1 vccd1 _16348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16279_ _16283_/CLK _16279_/D vssd1 vssd1 vccd1 vccd1 _16279_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07983_ _07983_/A _07983_/B vssd1 vssd1 vccd1 vccd1 _08177_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09722_ _15416_/Q _09727_/C _09490_/X vssd1 vssd1 vccd1 vccd1 _09724_/C sky130_fd_sc_hd__a21o_1
XFILLER_86_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09653_ _09652_/B _09652_/C _09596_/X vssd1 vssd1 vccd1 vccd1 _09654_/C sky130_fd_sc_hd__o21ai_1
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08604_ _09541_/A vssd1 vssd1 vccd1 vccd1 _08604_/X sky130_fd_sc_hd__clkbuf_2
X_09584_ _09643_/A _09584_/B _09588_/B vssd1 vssd1 vccd1 vccd1 _15392_/D sky130_fd_sc_hd__nor3_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08535_ _08535_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _08536_/B sky130_fd_sc_hd__nor2_1
XFILLER_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08466_ _08519_/A _08466_/B _08466_/C vssd1 vssd1 vccd1 vccd1 _08467_/A sky130_fd_sc_hd__and3_1
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08397_ _08397_/A _08397_/B vssd1 vssd1 vccd1 vccd1 _08397_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09018_ _09133_/A _09018_/B _09018_/C vssd1 vssd1 vccd1 vccd1 _09021_/B sky130_fd_sc_hd__or3_1
X_10290_ _10304_/C vssd1 vssd1 vccd1 vccd1 _10312_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13980_ _13980_/A _13980_/B _13985_/A vssd1 vssd1 vccd1 vccd1 _16099_/D sky130_fd_sc_hd__nor3_1
XFILLER_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12931_ _12962_/C vssd1 vssd1 vccd1 vccd1 _12968_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15650_ _15655_/CLK _15650_/D vssd1 vssd1 vccd1 vccd1 _15650_/Q sky130_fd_sc_hd__dfxtp_1
X_12862_ _15907_/Q _12861_/C _12631_/X vssd1 vssd1 vccd1 vccd1 _12863_/B sky130_fd_sc_hd__a21oi_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11813_ _15742_/Q _11814_/C _11812_/X vssd1 vssd1 vccd1 vccd1 _11813_/Y sky130_fd_sc_hd__a21oi_1
X_14601_ _14601_/A _14601_/B vssd1 vssd1 vccd1 vccd1 _14601_/X sky130_fd_sc_hd__or2_1
X_15581_ _15655_/CLK _15581_/D vssd1 vssd1 vccd1 vccd1 _15581_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _15895_/Q _12793_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12793_/Y sky130_fd_sc_hd__nand3_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14532_/A _14532_/B vssd1 vssd1 vccd1 vccd1 _14533_/B sky130_fd_sc_hd__and2_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11744_/A vssd1 vssd1 vccd1 vccd1 _15730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14466_/C vssd1 vssd1 vccd1 vccd1 _14474_/C sky130_fd_sc_hd__clkbuf_1
X_11675_ _11826_/A vssd1 vssd1 vccd1 vccd1 _11796_/A sky130_fd_sc_hd__clkbuf_2
X_16202_ _16204_/CLK _16202_/D vssd1 vssd1 vccd1 vccd1 _16202_/Q sky130_fd_sc_hd__dfxtp_1
X_13414_ _13412_/X _13410_/C _13413_/Y vssd1 vssd1 vccd1 vccd1 _15998_/D sky130_fd_sc_hd__a21oi_1
X_10626_ _10634_/B _10626_/B vssd1 vssd1 vccd1 vccd1 _10628_/A sky130_fd_sc_hd__or2_1
XFILLER_139_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14394_ _16186_/Q _14440_/B _14403_/C vssd1 vssd1 vccd1 vccd1 _14398_/A sky130_fd_sc_hd__and3_1
XFILLER_127_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16133_ _16222_/CLK _16133_/D vssd1 vssd1 vccd1 vccd1 _16133_/Q sky130_fd_sc_hd__dfxtp_1
X_13345_ _15987_/Q _13550_/B _13349_/C vssd1 vssd1 vccd1 vccd1 _13345_/Y sky130_fd_sc_hd__nand3_1
X_10557_ _10554_/X _10555_/Y _10556_/Y _10552_/C vssd1 vssd1 vccd1 vccd1 _10559_/B
+ sky130_fd_sc_hd__o211ai_1
X_16064_ _16148_/CLK _16064_/D vssd1 vssd1 vccd1 vccd1 _16064_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13276_ _15977_/Q _13484_/B _13276_/C vssd1 vssd1 vccd1 vccd1 _13276_/X sky130_fd_sc_hd__and3_1
X_10488_ _10503_/A _10488_/B _10488_/C vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__and3_1
XFILLER_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15015_ _14970_/X _15012_/A _15014_/X vssd1 vssd1 vccd1 vccd1 _15015_/Y sky130_fd_sc_hd__a21oi_1
X_12227_ _12227_/A vssd1 vssd1 vccd1 vccd1 _15805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12158_ _15796_/Q _12159_/C _12100_/X vssd1 vssd1 vccd1 vccd1 _12158_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11109_ _11110_/B _11110_/C _11110_/A vssd1 vssd1 vccd1 vccd1 _11111_/B sky130_fd_sc_hd__a21o_1
X_12089_ _12089_/A _12089_/B _12089_/C vssd1 vssd1 vccd1 vccd1 _12090_/C sky130_fd_sc_hd__nand3_1
XFILLER_111_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15917_ _15935_/CLK _15917_/D vssd1 vssd1 vccd1 vccd1 _15917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15848_ _15907_/CLK _15848_/D vssd1 vssd1 vccd1 vccd1 _15848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15779_ _15195_/Q _15779_/D vssd1 vssd1 vccd1 vccd1 _15779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08320_ _08359_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _08321_/B sky130_fd_sc_hd__xor2_2
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08251_ _08251_/A _08251_/B vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__xnor2_4
XFILLER_137_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08182_ _08182_/A _08043_/A vssd1 vssd1 vccd1 vccd1 _08182_/X sky130_fd_sc_hd__or2b_1
XFILLER_119_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07966_ _16197_/Q vssd1 vssd1 vccd1 vccd1 _14505_/C sky130_fd_sc_hd__inv_2
XFILLER_101_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09705_ _09760_/A _09708_/C vssd1 vssd1 vccd1 vccd1 _09705_/X sky130_fd_sc_hd__or2_1
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ _15458_/Q vssd1 vssd1 vccd1 vccd1 _10002_/A sky130_fd_sc_hd__clkinv_2
Xclkbuf_leaf_94_clk _15665_/CLK vssd1 vssd1 vccd1 vccd1 _15656_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09636_ _09636_/A vssd1 vssd1 vccd1 vccd1 _15400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09567_ _09565_/Y _09561_/C _09563_/X _09564_/Y vssd1 vssd1 vccd1 vccd1 _09568_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_130_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08518_ _08516_/Y _08508_/C _08512_/X _08514_/Y vssd1 vssd1 vccd1 vccd1 _08519_/C
+ sky130_fd_sc_hd__a211o_1
X_09498_ _15381_/Q _09508_/C _09497_/X vssd1 vssd1 vccd1 vccd1 _09498_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08449_ _08449_/A vssd1 vssd1 vccd1 vccd1 _15219_/D sky130_fd_sc_hd__clkbuf_1
X_11460_ _11454_/B _11455_/C _11457_/X _11458_/Y vssd1 vssd1 vccd1 vccd1 _11461_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_149_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10411_ _15521_/Q vssd1 vssd1 vccd1 vccd1 _10426_/C sky130_fd_sc_hd__inv_2
X_11391_ _11423_/C vssd1 vssd1 vccd1 vccd1 _11431_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13130_ _13130_/A vssd1 vssd1 vccd1 vccd1 _14261_/A sky130_fd_sc_hd__buf_2
XFILLER_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10342_ _10577_/A _10342_/B _10342_/C vssd1 vssd1 vccd1 vccd1 _10344_/B sky130_fd_sc_hd__or3_1
XFILLER_125_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _13059_/Y _13055_/C _13057_/X _13058_/Y vssd1 vssd1 vccd1 vccd1 _13062_/C
+ sky130_fd_sc_hd__a211o_1
X_10273_ _10271_/Y _10266_/C _10279_/A _10270_/Y vssd1 vssd1 vccd1 vccd1 _10279_/B
+ sky130_fd_sc_hd__a211oi_1
X_12012_ _12068_/A _12015_/C vssd1 vssd1 vccd1 vccd1 _12012_/X sky130_fd_sc_hd__or2_1
XFILLER_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13963_ _15186_/A _13963_/B vssd1 vssd1 vccd1 vccd1 _13964_/B sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_85_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15449_/CLK sky130_fd_sc_hd__clkbuf_16
X_15702_ _15794_/CLK _15702_/D vssd1 vssd1 vccd1 vccd1 _15702_/Q sky130_fd_sc_hd__dfxtp_2
X_12914_ _15916_/Q _13078_/B _12914_/C vssd1 vssd1 vccd1 vccd1 _12923_/B sky130_fd_sc_hd__and3_1
X_13894_ _16087_/Q _13903_/C _13893_/X vssd1 vssd1 vccd1 vccd1 _13896_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15633_ _15194_/Q _15633_/D vssd1 vssd1 vccd1 vccd1 _15633_/Q sky130_fd_sc_hd__dfxtp_1
X_12845_ _15905_/Q _12954_/B _12854_/C vssd1 vssd1 vccd1 vccd1 _12845_/X sky130_fd_sc_hd__and3_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15655_/CLK _15564_/D vssd1 vssd1 vccd1 vccd1 _15564_/Q sky130_fd_sc_hd__dfxtp_1
X_12776_ _12776_/A vssd1 vssd1 vccd1 vccd1 _15892_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11727_/A _11727_/B _11727_/C vssd1 vssd1 vccd1 vccd1 _11729_/B sky130_fd_sc_hd__or3_1
X_14515_ _14520_/A _14514_/Y _14510_/B _14511_/C vssd1 vssd1 vccd1 vccd1 _14517_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15495_ _15224_/Q _15495_/D vssd1 vssd1 vccd1 vccd1 _15495_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ _15716_/Q _11887_/B _11662_/C vssd1 vssd1 vccd1 vccd1 _11658_/Y sky130_fd_sc_hd__nand3_1
X_14446_ _14443_/B _14442_/Y _14443_/A vssd1 vssd1 vccd1 vccd1 _14446_/Y sky130_fd_sc_hd__o21bai_1
X_10609_ _15554_/Q _10609_/B _10617_/C vssd1 vssd1 vccd1 vccd1 _10609_/X sky130_fd_sc_hd__and3_1
XFILLER_127_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14377_ _14389_/C vssd1 vssd1 vccd1 vccd1 _14403_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11589_ _11589_/A vssd1 vssd1 vccd1 vccd1 _15705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13328_ _15986_/Q _13327_/C _13277_/X vssd1 vssd1 vccd1 vccd1 _13328_/Y sky130_fd_sc_hd__a21oi_1
X_16116_ _16142_/CLK _16116_/D vssd1 vssd1 vccd1 vccd1 _16116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16047_ _16050_/CLK _16047_/D vssd1 vssd1 vccd1 vccd1 _16047_/Q sky130_fd_sc_hd__dfxtp_1
X_13259_ _13154_/X _13257_/C _13206_/X vssd1 vssd1 vccd1 vccd1 _13259_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ _15872_/Q _07820_/B vssd1 vssd1 vccd1 vccd1 _07821_/B sky130_fd_sc_hd__or2_1
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07751_ _10058_/A _07751_/B vssd1 vssd1 vccd1 vccd1 _07752_/B sky130_fd_sc_hd__xnor2_4
XFILLER_38_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_76_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15348_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07682_ _13654_/A vssd1 vssd1 vccd1 vccd1 _14099_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09421_ _09458_/A _09421_/B _09421_/C vssd1 vssd1 vccd1 vccd1 _09422_/A sky130_fd_sc_hd__and3_1
XFILLER_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _09350_/Y _09345_/C _09357_/A _09349_/Y vssd1 vssd1 vccd1 vccd1 _09357_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_21_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08303_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08352_/A sky130_fd_sc_hd__xnor2_1
X_09283_ _15348_/Q _09451_/B _09290_/C vssd1 vssd1 vccd1 vccd1 _09283_/X sky130_fd_sc_hd__and3_1
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08234_ _08234_/A _08234_/B vssd1 vssd1 vccd1 vccd1 _08234_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08165_ _15208_/Q _08279_/A vssd1 vssd1 vccd1 vccd1 _08166_/B sky130_fd_sc_hd__nand2_1
X_08096_ _08096_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08097_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08998_ _08996_/Y _08992_/C _08994_/X _08995_/Y vssd1 vssd1 vccd1 vccd1 _08999_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_102_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07949_ _09543_/A _07949_/B vssd1 vssd1 vccd1 vccd1 _07949_/X sky130_fd_sc_hd__or2_1
XFILLER_56_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_67_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15282_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10960_ _10960_/A _10960_/B _10960_/C vssd1 vssd1 vccd1 vccd1 _10961_/A sky130_fd_sc_hd__and3_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _09635_/A _09619_/B _09619_/C vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__and3_1
XFILLER_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10891_ _10888_/X _10889_/Y _10890_/Y _10886_/C vssd1 vssd1 vccd1 vccd1 _10893_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12630_ _15871_/Q _12861_/B _12630_/C vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__and3_1
XFILLER_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12561_ _12847_/A vssd1 vssd1 vccd1 vccd1 _12793_/B sky130_fd_sc_hd__buf_2
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11512_ _12654_/A vssd1 vssd1 vccd1 vccd1 _11512_/X sky130_fd_sc_hd__clkbuf_2
X_14300_ _14300_/A vssd1 vssd1 vccd1 vccd1 _14300_/X sky130_fd_sc_hd__buf_2
X_15280_ _16352_/CLK _15280_/D vssd1 vssd1 vccd1 vccd1 _15280_/Q sky130_fd_sc_hd__dfxtp_2
X_12492_ _15849_/Q _12720_/B _12492_/C vssd1 vssd1 vccd1 vccd1 _12492_/X sky130_fd_sc_hd__and3_1
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14231_ _14227_/Y _14230_/X _14196_/X vssd1 vssd1 vccd1 vccd1 _14231_/Y sky130_fd_sc_hd__a21oi_1
X_11443_ _15691_/Q _15690_/Q _15689_/Q _11273_/X vssd1 vssd1 vccd1 vccd1 _15683_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_137_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14162_ _14208_/A _14162_/B _14168_/A vssd1 vssd1 vccd1 vccd1 _16135_/D sky130_fd_sc_hd__nor3_1
X_11374_ _15673_/Q _11431_/B _11374_/C vssd1 vssd1 vccd1 vccd1 _11382_/B sky130_fd_sc_hd__and3_1
XFILLER_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ _13105_/B _13106_/C _13109_/X _13111_/Y vssd1 vssd1 vccd1 vccd1 _13114_/C
+ sky130_fd_sc_hd__a211o_1
X_10325_ _15510_/Q _10446_/B _10325_/C vssd1 vssd1 vccd1 vccd1 _10336_/A sky130_fd_sc_hd__and3_1
XFILLER_125_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14093_ _16123_/Q _14093_/B _14093_/C vssd1 vssd1 vccd1 vccd1 _14102_/A sky130_fd_sc_hd__and3_1
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13077_/A _13044_/B _13048_/A vssd1 vssd1 vccd1 vccd1 _15937_/D sky130_fd_sc_hd__nor3_1
X_10256_ _15498_/Q _10492_/B _10256_/C vssd1 vssd1 vccd1 vccd1 _10256_/Y sky130_fd_sc_hd__nand3_1
XFILLER_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10187_ _10188_/B _10188_/C _10188_/A vssd1 vssd1 vccd1 vccd1 _10189_/B sky130_fd_sc_hd__a21o_1
XFILLER_79_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_58_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _16344_/CLK sky130_fd_sc_hd__clkbuf_16
X_14995_ hold6/X _14994_/C _14917_/X vssd1 vssd1 vccd1 vccd1 _14996_/B sky130_fd_sc_hd__a21oi_1
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13946_ _16095_/Q _13945_/C _14088_/B vssd1 vssd1 vccd1 vccd1 _13946_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13877_ _16085_/Q _13981_/B _13885_/C vssd1 vssd1 vccd1 vccd1 _13881_/B sky130_fd_sc_hd__nand3_1
XFILLER_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _15194_/Q _15616_/D vssd1 vssd1 vccd1 vccd1 _15616_/Q sky130_fd_sc_hd__dfxtp_1
X_12828_ _12829_/B _12829_/C _12829_/A vssd1 vssd1 vccd1 vccd1 _12830_/B sky130_fd_sc_hd__a21o_1
XFILLER_62_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15547_ _15655_/CLK _15547_/D vssd1 vssd1 vccd1 vccd1 _15547_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12757_/B _12757_/C _12758_/X vssd1 vssd1 vccd1 vccd1 _12760_/C sky130_fd_sc_hd__o21ai_1
XFILLER_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15478_ _15483_/CLK _15478_/D vssd1 vssd1 vccd1 vccd1 _15478_/Q sky130_fd_sc_hd__dfxtp_1
X_14429_ _16193_/Q _14435_/C _14250_/X vssd1 vssd1 vccd1 vccd1 _14431_/C sky130_fd_sc_hd__a21o_1
XFILLER_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09970_ _09977_/A _09970_/B _09970_/C vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__and3_1
XFILLER_131_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08921_ _15292_/Q _08931_/C _08920_/X vssd1 vssd1 vccd1 vccd1 _08921_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08852_ _08909_/A _08852_/B _08856_/A vssd1 vssd1 vccd1 vccd1 _15280_/D sky130_fd_sc_hd__nor3_1
XFILLER_85_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07803_ _15809_/Q _15827_/Q vssd1 vssd1 vccd1 vccd1 _08049_/B sky130_fd_sc_hd__xor2_2
XFILLER_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08783_ _08839_/A _08783_/B _08783_/C vssd1 vssd1 vccd1 vccd1 _08785_/B sky130_fd_sc_hd__or3_1
XFILLER_69_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16273_/CLK sky130_fd_sc_hd__clkbuf_16
X_07734_ _15351_/Q _07734_/B vssd1 vssd1 vccd1 vccd1 _07735_/B sky130_fd_sc_hd__xnor2_2
XFILLER_84_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07665_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07667_/A sky130_fd_sc_hd__or2_1
X_09404_ _09693_/A vssd1 vssd1 vccd1 vccd1 _09404_/X sky130_fd_sc_hd__buf_2
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _09332_/X _09333_/Y _09334_/Y _09330_/C vssd1 vssd1 vccd1 vccd1 _09337_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09266_ _09266_/A _09266_/B _09266_/C vssd1 vssd1 vccd1 vccd1 _09267_/C sky130_fd_sc_hd__nand3_1
Xclkbuf_opt_1_0_clk _15665_/CLK vssd1 vssd1 vccd1 vccd1 _15692_/CLK sky130_fd_sc_hd__clkbuf_16
X_08217_ _08217_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08218_/B sky130_fd_sc_hd__and2_1
X_09197_ _09211_/C vssd1 vssd1 vccd1 vccd1 _09222_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_08148_ _15368_/Q _08148_/B vssd1 vssd1 vccd1 vccd1 _08148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08079_ _08222_/A _08222_/B vssd1 vssd1 vccd1 vccd1 _08080_/B sky130_fd_sc_hd__xor2_1
XFILLER_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10110_ _10110_/A vssd1 vssd1 vccd1 vccd1 _10338_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11090_ _11090_/A _11090_/B vssd1 vssd1 vccd1 vccd1 _11094_/C sky130_fd_sc_hd__nor2_1
XFILLER_96_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10041_ _10039_/Y _10035_/C _10047_/A _10038_/Y vssd1 vssd1 vccd1 vccd1 _10047_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_121_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13800_ _16069_/Q _13805_/C _13598_/X vssd1 vssd1 vccd1 vccd1 _13800_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_75_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11992_ _15770_/Q _12000_/C _11760_/X vssd1 vssd1 vccd1 vccd1 _11992_/Y sky130_fd_sc_hd__a21oi_1
X_14780_ _14979_/A vssd1 vssd1 vccd1 vccd1 _14946_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13731_ _16057_/Q _14074_/B _13738_/C vssd1 vssd1 vccd1 vccd1 _13734_/B sky130_fd_sc_hd__nand3_1
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10943_ _10936_/B _10937_/C _10939_/X _10941_/Y vssd1 vssd1 vccd1 vccd1 _10944_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 _15665_/CLK sky130_fd_sc_hd__clkbuf_2
X_10874_ _15595_/Q _11161_/B _10882_/C vssd1 vssd1 vccd1 vccd1 _10879_/A sky130_fd_sc_hd__and3_1
X_13662_ _13662_/A _13662_/B _13662_/C vssd1 vssd1 vccd1 vccd1 _13664_/B sky130_fd_sc_hd__or3_1
XFILLER_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15401_ _15484_/CLK _15401_/D vssd1 vssd1 vccd1 vccd1 _15401_/Q sky130_fd_sc_hd__dfxtp_1
X_12613_ _12621_/A _12613_/B _12613_/C vssd1 vssd1 vccd1 vccd1 _12614_/A sky130_fd_sc_hd__and3_1
X_13593_ _13589_/X _13590_/Y _13592_/Y _13587_/C vssd1 vssd1 vccd1 vccd1 _13595_/B
+ sky130_fd_sc_hd__o211ai_1
X_15332_ _15339_/CLK _15332_/D vssd1 vssd1 vccd1 vccd1 _15332_/Q sky130_fd_sc_hd__dfxtp_1
X_12544_ _12565_/A _12544_/B _12544_/C vssd1 vssd1 vccd1 vccd1 _12545_/A sky130_fd_sc_hd__and3_1
XFILLER_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15263_ _15274_/CLK _15263_/D vssd1 vssd1 vccd1 vccd1 _15263_/Q sky130_fd_sc_hd__dfxtp_1
X_12475_ _12475_/A vssd1 vssd1 vccd1 vccd1 _15844_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14214_ _14214_/A vssd1 vssd1 vccd1 vccd1 _16145_/D sky130_fd_sc_hd__clkbuf_1
X_11426_ _15681_/Q _11431_/C _11425_/X vssd1 vssd1 vccd1 vccd1 _11426_/Y sky130_fd_sc_hd__a21oi_1
X_15194_ _15224_/Q _15194_/D vssd1 vssd1 vccd1 vccd1 _15194_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_6 _15176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14145_ _14320_/A _14145_/B vssd1 vssd1 vccd1 vccd1 _14146_/B sky130_fd_sc_hd__and2_1
X_11357_ _11355_/Y _11351_/C _11353_/X _11354_/Y vssd1 vssd1 vccd1 vccd1 _11358_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10308_ _10323_/A _10308_/B _10308_/C vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__and3_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14076_ _14077_/B _14077_/C _14077_/A vssd1 vssd1 vccd1 vccd1 _14078_/B sky130_fd_sc_hd__a21o_1
X_11288_ _11288_/A vssd1 vssd1 vccd1 vccd1 _15658_/D sky130_fd_sc_hd__clkbuf_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _13199_/A _13031_/C vssd1 vssd1 vccd1 vccd1 _13027_/X sky130_fd_sc_hd__or2_1
X_10239_ _15496_/Q _10239_/B _10247_/C vssd1 vssd1 vccd1 vccd1 _10244_/A sky130_fd_sc_hd__and3_1
XFILLER_94_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14978_ _15023_/A _14978_/B _14984_/A vssd1 vssd1 vccd1 vccd1 _16315_/D sky130_fd_sc_hd__nor3_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13929_ _14372_/A vssd1 vssd1 vccd1 vccd1 _15013_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09120_ _15321_/Q _09238_/B _09125_/C vssd1 vssd1 vccd1 vccd1 _09120_/Y sky130_fd_sc_hd__nand3_1
X_09051_ _09051_/A vssd1 vssd1 vccd1 vccd1 _15310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08002_ _08002_/A _08188_/A vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__xnor2_4
XFILLER_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09953_ _15452_/Q _09958_/C _09778_/X vssd1 vssd1 vccd1 vccd1 _09955_/C sky130_fd_sc_hd__a21o_1
XFILLER_103_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08904_ _08919_/C vssd1 vssd1 vccd1 vccd1 _08931_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09884_ _10751_/A vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__clkbuf_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _08835_/A _08835_/B vssd1 vssd1 vccd1 vccd1 _08839_/C sky130_fd_sc_hd__nor2_1
XFILLER_85_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08766_ _08766_/A vssd1 vssd1 vccd1 vccd1 _15266_/D sky130_fd_sc_hd__clkbuf_1
X_07717_ _15566_/Q vssd1 vssd1 vccd1 vccd1 _10700_/A sky130_fd_sc_hd__clkinv_4
X_08697_ _08704_/A _08697_/B _08697_/C vssd1 vssd1 vccd1 vccd1 _08698_/A sky130_fd_sc_hd__and3_1
XFILLER_14_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07648_ _10950_/C vssd1 vssd1 vccd1 vccd1 _15171_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09318_ _15353_/Q _09372_/B _09326_/C vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__and3_1
XFILLER_139_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10590_ _15551_/Q _10590_/B _10596_/C vssd1 vssd1 vccd1 vccd1 _10593_/B sky130_fd_sc_hd__nand3_1
X_09249_ _09247_/A _09247_/B _09248_/X vssd1 vssd1 vccd1 vccd1 _15340_/D sky130_fd_sc_hd__a21oi_1
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12260_ _12281_/A _12260_/B _12260_/C vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__and3_1
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11211_ _11211_/A vssd1 vssd1 vccd1 vccd1 _15646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12191_ _12191_/A vssd1 vssd1 vccd1 vccd1 _15799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11142_ _11220_/A _11142_/B _11146_/B vssd1 vssd1 vccd1 vccd1 _15635_/D sky130_fd_sc_hd__nor3_1
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11073_ _15625_/Q _11073_/B _11078_/C vssd1 vssd1 vccd1 vccd1 _11073_/Y sky130_fd_sc_hd__nand3_1
X_15950_ _15956_/CLK _15950_/D vssd1 vssd1 vccd1 vccd1 _15950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10024_ _15462_/Q _10199_/B _10024_/C vssd1 vssd1 vccd1 vccd1 _10024_/Y sky130_fd_sc_hd__nand3_1
X_14901_ _14901_/A vssd1 vssd1 vccd1 vccd1 _14901_/X sky130_fd_sc_hd__buf_2
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15881_ _15961_/CLK _15881_/D vssd1 vssd1 vccd1 vccd1 _15881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14832_ _14936_/A vssd1 vssd1 vccd1 vccd1 _14915_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14763_ _14847_/A _14769_/C vssd1 vssd1 vccd1 vccd1 _14763_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11975_ _11975_/A _11975_/B _11975_/C vssd1 vssd1 vccd1 vccd1 _11976_/C sky130_fd_sc_hd__nand3_1
XFILLER_32_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13714_ _13712_/A _13712_/B _13713_/X vssd1 vssd1 vccd1 vccd1 _16050_/D sky130_fd_sc_hd__a21oi_1
X_10926_ _10939_/B vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14694_ _14892_/A vssd1 vssd1 vccd1 vccd1 _14694_/X sky130_fd_sc_hd__clkbuf_2
X_13645_ _13643_/Y _13638_/C _13641_/X _13642_/Y vssd1 vssd1 vccd1 vccd1 _13646_/C
+ sky130_fd_sc_hd__a211o_1
X_10857_ _10863_/B _10857_/B vssd1 vssd1 vccd1 vccd1 _10859_/A sky130_fd_sc_hd__or2_1
XFILLER_13_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _16364_/CLK _16364_/D vssd1 vssd1 vccd1 vccd1 _16364_/Q sky130_fd_sc_hd__dfxtp_1
X_13576_ _13604_/A _13576_/B _13580_/A vssd1 vssd1 vccd1 vccd1 _16027_/D sky130_fd_sc_hd__nor3_1
XFILLER_13_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ _10786_/Y _10781_/C _10783_/X _10784_/Y vssd1 vssd1 vccd1 vccd1 _10789_/C
+ sky130_fd_sc_hd__a211o_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15315_ _15333_/CLK _15315_/D vssd1 vssd1 vccd1 vccd1 _15315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12527_ _12583_/A _12527_/B _12527_/C vssd1 vssd1 vccd1 vccd1 _12529_/B sky130_fd_sc_hd__or3_1
X_16295_ _16321_/CLK _16295_/D vssd1 vssd1 vccd1 vccd1 _16295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15246_ _15254_/CLK _15246_/D vssd1 vssd1 vccd1 vccd1 _15246_/Q sky130_fd_sc_hd__dfxtp_1
X_12458_ _15842_/Q _12458_/B _12462_/C vssd1 vssd1 vccd1 vccd1 _12458_/Y sky130_fd_sc_hd__nand3_1
XFILLER_126_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11409_ _15678_/Q _11409_/B _11409_/C vssd1 vssd1 vccd1 vccd1 _11409_/Y sky130_fd_sc_hd__nand3_1
XFILLER_141_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12389_ _12396_/A _12389_/B _12389_/C vssd1 vssd1 vccd1 vccd1 _12390_/A sky130_fd_sc_hd__and3_1
X_15177_ _16367_/Q _15176_/C _13950_/B vssd1 vssd1 vccd1 vccd1 _15178_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14128_ _14122_/B _14123_/C _14132_/A _14126_/Y vssd1 vssd1 vccd1 vccd1 _14132_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14059_ _14326_/A vssd1 vssd1 vccd1 vccd1 _14059_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ _08648_/A _08620_/B _08620_/C vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__and3_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _13043_/B vssd1 vssd1 vccd1 vccd1 _08794_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08482_ _08611_/A hold2/X _08488_/A vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__nor3_1
XFILLER_63_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09103_ _15320_/Q _09105_/C _08929_/X vssd1 vssd1 vccd1 vccd1 _09103_/Y sky130_fd_sc_hd__a21oi_1
X_09034_ _15309_/Q _09039_/C _08913_/X vssd1 vssd1 vccd1 vccd1 _09036_/C sky130_fd_sc_hd__a21o_1
XFILLER_136_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09936_ _10049_/A _09939_/C vssd1 vssd1 vccd1 vccd1 _09936_/X sky130_fd_sc_hd__or2_1
XFILLER_132_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09867_ _15438_/Q _09867_/B _09867_/C vssd1 vssd1 vccd1 vccd1 _09877_/A sky130_fd_sc_hd__and3_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _15275_/Q _08996_/B _08823_/C vssd1 vssd1 vccd1 vccd1 _08818_/Y sky130_fd_sc_hd__nand3_1
XFILLER_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09798_ _09796_/Y _09790_/C _09793_/X _09795_/Y vssd1 vssd1 vccd1 vccd1 _09799_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _08765_/A _08749_/B _08749_/C vssd1 vssd1 vccd1 vccd1 _08750_/A sky130_fd_sc_hd__and3_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11760_ _12048_/A vssd1 vssd1 vccd1 vccd1 _11760_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10732_/A _10711_/B _10711_/C vssd1 vssd1 vccd1 vccd1 _10712_/A sky130_fd_sc_hd__and3_1
XFILLER_26_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11689_/X _11690_/Y _11686_/B _11687_/C vssd1 vssd1 vccd1 vccd1 _11693_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10642_ _10679_/C vssd1 vssd1 vccd1 vccd1 _10685_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13430_ _16004_/Q _13484_/B _13430_/C vssd1 vssd1 vccd1 vccd1 _13430_/X sky130_fd_sc_hd__and3_1
XFILLER_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13361_ _13361_/A vssd1 vssd1 vccd1 vccd1 _15988_/D sky130_fd_sc_hd__clkbuf_1
X_10573_ _10573_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _10577_/C sky130_fd_sc_hd__nor2_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15100_ _15135_/A _15100_/B _15100_/C vssd1 vssd1 vccd1 vccd1 _15101_/A sky130_fd_sc_hd__and3_1
X_12312_ _15821_/Q _12317_/C _12086_/X vssd1 vssd1 vccd1 vccd1 _12314_/C sky130_fd_sc_hd__a21o_1
XFILLER_139_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16080_ _16103_/CLK _16080_/D vssd1 vssd1 vccd1 vccd1 _16080_/Q sky130_fd_sc_hd__dfxtp_1
X_13292_ _15979_/Q _13297_/C _14605_/B vssd1 vssd1 vccd1 vccd1 _13292_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12243_ _12299_/A _12243_/B _12243_/C vssd1 vssd1 vccd1 vccd1 _12245_/B sky130_fd_sc_hd__or3_1
X_15031_ _16330_/Q _15031_/B _15036_/C vssd1 vssd1 vccd1 vccd1 _15039_/A sky130_fd_sc_hd__and3_1
X_12174_ _15797_/Q _12174_/B _12178_/C vssd1 vssd1 vccd1 vccd1 _12174_/Y sky130_fd_sc_hd__nand3_1
XFILLER_123_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11125_ _11125_/A vssd1 vssd1 vccd1 vccd1 _15633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11056_ _11056_/A vssd1 vssd1 vccd1 vccd1 _15622_/D sky130_fd_sc_hd__clkbuf_1
X_15933_ _15196_/Q _15933_/D vssd1 vssd1 vccd1 vccd1 _15933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10007_ _10007_/A vssd1 vssd1 vccd1 vccd1 _10239_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15864_ _07603_/A _15864_/D vssd1 vssd1 vccd1 vccd1 _15864_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14815_ _15014_/A vssd1 vssd1 vccd1 vccd1 _14815_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15795_ _15195_/Q _15795_/D vssd1 vssd1 vccd1 vccd1 _15795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14746_ _14747_/B _14747_/C _14747_/A vssd1 vssd1 vccd1 vccd1 _14748_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11958_ _12015_/A _11958_/B _11958_/C vssd1 vssd1 vccd1 vccd1 _11960_/B sky130_fd_sc_hd__or3_1
XFILLER_60_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10909_ _10931_/A _10909_/B _10914_/B vssd1 vssd1 vccd1 vccd1 _15599_/D sky130_fd_sc_hd__nor3_1
X_14677_ _16250_/Q _14755_/B _14677_/C vssd1 vssd1 vccd1 vccd1 _14679_/A sky130_fd_sc_hd__and3_1
X_11889_ _11887_/Y _11883_/C _11894_/A _11886_/Y vssd1 vssd1 vccd1 vccd1 _11894_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13628_ _16039_/Q _13628_/B _13634_/C vssd1 vssd1 vccd1 vccd1 _13631_/B sky130_fd_sc_hd__nand3_1
XFILLER_20_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16347_ _16364_/CLK _16347_/D vssd1 vssd1 vccd1 vccd1 _16347_/Q sky130_fd_sc_hd__dfxtp_1
X_13559_ _13713_/A _13561_/C vssd1 vssd1 vccd1 vccd1 _13559_/X sky130_fd_sc_hd__or2_1
XFILLER_146_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16278_ _16317_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _16278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15229_ _15926_/CLK _15229_/D vssd1 vssd1 vccd1 vccd1 _15229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07982_ _08180_/A _08180_/B vssd1 vssd1 vccd1 vccd1 _07983_/B sky130_fd_sc_hd__xor2_2
XFILLER_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09721_ _15416_/Q _09721_/B _09727_/C vssd1 vssd1 vccd1 vccd1 _09724_/B sky130_fd_sc_hd__nand3_1
XFILLER_68_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09652_ _09708_/A _09652_/B _09652_/C vssd1 vssd1 vccd1 vccd1 _09654_/B sky130_fd_sc_hd__or3_1
XFILLER_95_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08603_ _08603_/A vssd1 vssd1 vccd1 vccd1 _15242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09583_ _09581_/Y _09575_/C _09588_/A _09578_/Y vssd1 vssd1 vccd1 vccd1 _09588_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_103_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ _08540_/B _08534_/B vssd1 vssd1 vccd1 vccd1 _08536_/A sky130_fd_sc_hd__or2_1
X_08465_ _08465_/A _08465_/B _08465_/C vssd1 vssd1 vccd1 vccd1 _08466_/C sky130_fd_sc_hd__or3_1
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08396_ _08403_/B _08452_/B vssd1 vssd1 vccd1 vccd1 _08397_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09017_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09058_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09919_ _15445_/Q _10150_/B _09925_/C vssd1 vssd1 vccd1 vccd1 _09919_/Y sky130_fd_sc_hd__nand3_1
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12930_ _12949_/C vssd1 vssd1 vccd1 vccd1 _12962_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12861_ _15907_/Q _12861_/B _12861_/C vssd1 vssd1 vccd1 vccd1 _12869_/B sky130_fd_sc_hd__and3_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14600_/A _14600_/B vssd1 vssd1 vccd1 vccd1 _14600_/Y sky130_fd_sc_hd__nor2_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _12100_/A vssd1 vssd1 vccd1 vccd1 _11812_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _15194_/Q _15580_/D vssd1 vssd1 vccd1 vccd1 _15580_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _15896_/Q _12798_/C _12616_/X vssd1 vssd1 vccd1 vccd1 _12792_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14524_/Y _14525_/X _14527_/B vssd1 vssd1 vccd1 vccd1 _14532_/B sky130_fd_sc_hd__o21a_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11743_ _11765_/A _11743_/B _11743_/C vssd1 vssd1 vccd1 vccd1 _11744_/A sky130_fd_sc_hd__and3_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _16214_/Q _16213_/Q _16212_/Q _14421_/X vssd1 vssd1 vccd1 vccd1 _16197_/D
+ sky130_fd_sc_hd__o31a_1
X_11674_ _15727_/Q _15726_/Q _15725_/Q _11560_/X vssd1 vssd1 vccd1 vccd1 _15719_/D
+ sky130_fd_sc_hd__o31a_1
X_16201_ _16204_/CLK _16201_/D vssd1 vssd1 vccd1 vccd1 _16201_/Q sky130_fd_sc_hd__dfxtp_1
X_13413_ _13362_/X _13410_/C _13206_/X vssd1 vssd1 vccd1 vccd1 _13413_/Y sky130_fd_sc_hd__o21ai_1
X_10625_ _15556_/Q _10623_/C _10624_/X vssd1 vssd1 vccd1 vccd1 _10626_/B sky130_fd_sc_hd__a21oi_1
X_14393_ _14427_/A _14393_/B _14397_/B vssd1 vssd1 vccd1 vccd1 _16182_/D sky130_fd_sc_hd__nor3_1
XFILLER_128_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16132_ _16222_/CLK _16132_/D vssd1 vssd1 vccd1 vccd1 _16132_/Q sky130_fd_sc_hd__dfxtp_1
X_10556_ _15544_/Q _10729_/B _10561_/C vssd1 vssd1 vccd1 vccd1 _10556_/Y sky130_fd_sc_hd__nand3_1
X_13344_ _14395_/A vssd1 vssd1 vccd1 vccd1 _13550_/B sky130_fd_sc_hd__buf_2
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ _16148_/CLK _16063_/D vssd1 vssd1 vccd1 vccd1 _16063_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10487_ _10481_/B _10482_/C _10484_/X _10485_/Y vssd1 vssd1 vccd1 vccd1 _10488_/C
+ sky130_fd_sc_hd__a211o_1
X_13275_ _13275_/A vssd1 vssd1 vccd1 vccd1 _13484_/B sky130_fd_sc_hd__buf_2
XFILLER_108_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15014_ _15014_/A vssd1 vssd1 vccd1 vccd1 _15014_/X sky130_fd_sc_hd__clkbuf_2
X_12226_ _12226_/A _12226_/B _12226_/C vssd1 vssd1 vccd1 vccd1 _12227_/A sky130_fd_sc_hd__and3_1
XFILLER_123_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12157_ _15796_/Q _12383_/B _12159_/C vssd1 vssd1 vccd1 vccd1 _12157_/X sky130_fd_sc_hd__and3_1
XFILLER_78_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _15632_/Q _11113_/C _10933_/X vssd1 vssd1 vccd1 vccd1 _11110_/C sky130_fd_sc_hd__a21o_1
XFILLER_111_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12088_ _12089_/B _12089_/C _12089_/A vssd1 vssd1 vccd1 vccd1 _12090_/B sky130_fd_sc_hd__a21o_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11039_ _11036_/B _11036_/C _11038_/X vssd1 vssd1 vccd1 vccd1 _11040_/C sky130_fd_sc_hd__o21ai_1
X_15916_ _15196_/Q _15916_/D vssd1 vssd1 vccd1 vccd1 _15916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15847_ _15907_/CLK _15847_/D vssd1 vssd1 vccd1 vccd1 _15847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15778_ _15794_/CLK _15778_/D vssd1 vssd1 vccd1 vccd1 _15778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14729_ _07688_/X _14731_/C _14695_/X vssd1 vssd1 vccd1 vccd1 _14730_/B sky130_fd_sc_hd__o21ai_1
X_08250_ _08250_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08251_/B sky130_fd_sc_hd__nor2_2
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08181_ _07983_/A _07983_/B _08180_/Y vssd1 vssd1 vccd1 vccd1 _08200_/A sky130_fd_sc_hd__a21o_1
XFILLER_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07965_ _16179_/Q vssd1 vssd1 vccd1 vccd1 _14426_/C sky130_fd_sc_hd__clkinv_2
X_09704_ _09704_/A _09704_/B vssd1 vssd1 vccd1 vccd1 _09708_/C sky130_fd_sc_hd__nor2_1
XFILLER_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07896_ _15386_/Q vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__clkinv_2
XFILLER_67_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09635_ _09635_/A _09635_/B _09635_/C vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__and3_1
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09566_ _09563_/X _09564_/Y _09565_/Y _09561_/C vssd1 vssd1 vccd1 vccd1 _09568_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08517_ _08512_/X _08514_/Y _08516_/Y _08508_/C vssd1 vssd1 vccd1 vccd1 _08519_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09497_ _13051_/B vssd1 vssd1 vccd1 vccd1 _09497_/X sky130_fd_sc_hd__buf_2
X_08448_ _08448_/A _08448_/B vssd1 vssd1 vccd1 vccd1 _08449_/A sky130_fd_sc_hd__and2_1
XFILLER_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _08379_/A vssd1 vssd1 vccd1 vccd1 _15210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10410_ _15529_/Q _15528_/Q _15527_/Q _10409_/X vssd1 vssd1 vccd1 vccd1 _15521_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ _11409_/C vssd1 vssd1 vccd1 vccd1 _11423_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ _10341_/A vssd1 vssd1 vccd1 vccd1 _10577_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ _13057_/X _13058_/Y _13059_/Y _13055_/C vssd1 vssd1 vccd1 vccd1 _13062_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10272_ _10279_/A _10270_/Y _10271_/Y _10266_/C vssd1 vssd1 vccd1 vccd1 _10274_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12011_ _12011_/A _12011_/B vssd1 vssd1 vccd1 vccd1 _12015_/C sky130_fd_sc_hd__nor2_1
XFILLER_133_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13962_ _13956_/Y _13957_/X _13959_/B vssd1 vssd1 vccd1 vccd1 _13963_/B sky130_fd_sc_hd__o21a_1
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15701_ _15701_/CLK _15701_/D vssd1 vssd1 vccd1 vccd1 _15701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12913_ _12934_/A _12913_/B _12917_/B vssd1 vssd1 vccd1 vccd1 _15914_/D sky130_fd_sc_hd__nor3_1
XFILLER_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13893_ _14598_/B vssd1 vssd1 vccd1 vccd1 _13893_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15632_ _15194_/Q _15632_/D vssd1 vssd1 vccd1 vccd1 _15632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12844_ _12844_/A vssd1 vssd1 vccd1 vccd1 _15903_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15655_/CLK _15563_/D vssd1 vssd1 vccd1 vccd1 _15563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12775_ _12796_/A _12775_/B _12775_/C vssd1 vssd1 vccd1 vccd1 _12776_/A sky130_fd_sc_hd__and3_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _16212_/Q _14513_/C _14634_/B vssd1 vssd1 vccd1 vccd1 _14514_/Y sky130_fd_sc_hd__a21oi_1
X_11726_ _11842_/A vssd1 vssd1 vccd1 vccd1 _11765_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15512_/CLK _15494_/D vssd1 vssd1 vccd1 vccd1 _15494_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14445_ _14443_/A _14443_/B _14442_/Y _14444_/Y vssd1 vssd1 vccd1 vccd1 _16192_/D
+ sky130_fd_sc_hd__o31a_1
X_11657_ _12230_/A vssd1 vssd1 vccd1 vccd1 _11887_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ _10608_/A vssd1 vssd1 vccd1 vccd1 _15552_/D sky130_fd_sc_hd__clkbuf_1
X_14376_ _14380_/C vssd1 vssd1 vccd1 vccd1 _14389_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11588_ _11597_/A _11588_/B _11588_/C vssd1 vssd1 vccd1 vccd1 _11589_/A sky130_fd_sc_hd__and3_1
XFILLER_128_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16115_ _16222_/CLK _16115_/D vssd1 vssd1 vccd1 vccd1 _16115_/Q sky130_fd_sc_hd__dfxtp_1
X_13327_ _15986_/Q _13484_/B _13327_/C vssd1 vssd1 vccd1 vccd1 _13327_/X sky130_fd_sc_hd__and3_1
XFILLER_143_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10539_ _10539_/A vssd1 vssd1 vccd1 vccd1 _15541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _16060_/CLK _16046_/D vssd1 vssd1 vccd1 vccd1 _16046_/Q sky130_fd_sc_hd__dfxtp_2
X_13258_ _13258_/A vssd1 vssd1 vccd1 vccd1 _15970_/D sky130_fd_sc_hd__clkbuf_1
X_12209_ _15804_/Q _12216_/C _12093_/X vssd1 vssd1 vccd1 vccd1 _12209_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13189_ _15960_/Q _13293_/B _13193_/C vssd1 vssd1 vccd1 vccd1 _13189_/Y sky130_fd_sc_hd__nand3_1
XFILLER_111_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07750_ _07750_/A _07750_/B vssd1 vssd1 vccd1 vccd1 _07751_/B sky130_fd_sc_hd__nand2_2
XFILLER_84_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07681_ _11424_/A vssd1 vssd1 vccd1 vccd1 _13654_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09420_ _09419_/B _09419_/C _09307_/X vssd1 vssd1 vccd1 vccd1 _09421_/C sky130_fd_sc_hd__o21ai_1
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ _09357_/A _09349_/Y _09350_/Y _09345_/C vssd1 vssd1 vccd1 vccd1 _09353_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08302_ _08211_/A _08062_/A _08062_/B _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1
+ _08351_/B sky130_fd_sc_hd__o32a_2
X_09282_ _09282_/A vssd1 vssd1 vccd1 vccd1 _15346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08233_ _08300_/B _08233_/B vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__xnor2_4
XFILLER_21_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08164_ spike_out[1] vssd1 vssd1 vccd1 vccd1 _08279_/A sky130_fd_sc_hd__inv_2
XFILLER_118_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08095_ _08096_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08238_/A sky130_fd_sc_hd__or2_2
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08997_ _08994_/X _08995_/Y _08996_/Y _08992_/C vssd1 vssd1 vccd1 vccd1 _08999_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07948_ _09196_/A _07934_/B _07933_/B vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__o21ai_4
XFILLER_68_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07879_ _07879_/A _07879_/B vssd1 vssd1 vccd1 vccd1 _07880_/B sky130_fd_sc_hd__nand2_2
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09618_ _09612_/B _09613_/C _09615_/X _09616_/Y vssd1 vssd1 vccd1 vccd1 _09619_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10890_ _15597_/Q _11121_/B _10890_/C vssd1 vssd1 vccd1 vccd1 _10890_/Y sky130_fd_sc_hd__nand3_1
X_09549_ _09643_/A _09549_/B _09553_/A vssd1 vssd1 vccd1 vccd1 _15387_/D sky130_fd_sc_hd__nor3_1
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12560_ _15860_/Q _12568_/C _12332_/X vssd1 vssd1 vccd1 vccd1 _12560_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11511_ input2/X vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__buf_4
XFILLER_12_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12491_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12720_/B sky130_fd_sc_hd__buf_2
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14230_ _14228_/X _14230_/B vssd1 vssd1 vccd1 vccd1 _14230_/X sky130_fd_sc_hd__and2b_1
X_11442_ _11442_/A vssd1 vssd1 vccd1 vccd1 _15682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11373_ _11373_/A _11373_/B _11377_/B vssd1 vssd1 vccd1 vccd1 _15671_/D sky130_fd_sc_hd__nor3_1
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14161_ _16138_/Q _14337_/B _14161_/C vssd1 vssd1 vccd1 vccd1 _14168_/A sky130_fd_sc_hd__and3_1
X_10324_ _10324_/A vssd1 vssd1 vccd1 vccd1 _15508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13112_ _13109_/X _13111_/Y _13105_/B _13106_/C vssd1 vssd1 vccd1 vccd1 _13114_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_125_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14092_ _14092_/A vssd1 vssd1 vccd1 vccd1 _16120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10255_ _10548_/A vssd1 vssd1 vccd1 vccd1 _10492_/B sky130_fd_sc_hd__buf_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _15938_/Q _13043_/B _13051_/C vssd1 vssd1 vccd1 vccd1 _13048_/A sky130_fd_sc_hd__and3_1
XFILLER_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10186_ _15488_/Q _10191_/C _10068_/X vssd1 vssd1 vccd1 vccd1 _10188_/C sky130_fd_sc_hd__a21o_1
XFILLER_78_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14994_ hold6/X _15142_/B _14994_/C vssd1 vssd1 vccd1 vccd1 _14996_/A sky130_fd_sc_hd__and3_1
XFILLER_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13945_ _16095_/Q _14988_/A _13945_/C vssd1 vssd1 vccd1 vccd1 _13952_/A sky130_fd_sc_hd__and3_1
XFILLER_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13876_ _14291_/A vssd1 vssd1 vccd1 vccd1 _13981_/B sky130_fd_sc_hd__buf_2
XFILLER_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15615_ _15194_/Q _15615_/D vssd1 vssd1 vccd1 vccd1 _15615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12827_ _15902_/Q _12832_/C _12654_/X vssd1 vssd1 vccd1 vccd1 _12829_/C sky130_fd_sc_hd__a21o_1
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15546_ _15655_/CLK _15546_/D vssd1 vssd1 vccd1 vccd1 _15546_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12758_/A vssd1 vssd1 vccd1 vccd1 _12758_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _11709_/A vssd1 vssd1 vccd1 vccd1 _15724_/D sky130_fd_sc_hd__clkbuf_1
X_15477_ _15483_/CLK _15477_/D vssd1 vssd1 vccd1 vccd1 _15477_/Q sky130_fd_sc_hd__dfxtp_2
X_12689_ _12804_/A _12689_/B _12693_/B vssd1 vssd1 vccd1 vccd1 _15878_/D sky130_fd_sc_hd__nor3_1
XFILLER_147_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14428_ _16193_/Q _14468_/B _14435_/C vssd1 vssd1 vccd1 vccd1 _14431_/B sky130_fd_sc_hd__nand3_1
XFILLER_128_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14359_ _14357_/X _14359_/B vssd1 vssd1 vccd1 vccd1 _14359_/X sky130_fd_sc_hd__and2b_1
XFILLER_115_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16029_ _16040_/CLK _16029_/D vssd1 vssd1 vccd1 vccd1 _16029_/Q sky130_fd_sc_hd__dfxtp_1
X_08920_ _13051_/B vssd1 vssd1 vccd1 vccd1 _08920_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08851_ _15281_/Q _09088_/B _08859_/C vssd1 vssd1 vccd1 vccd1 _08856_/A sky130_fd_sc_hd__and3_1
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07802_ _16170_/Q vssd1 vssd1 vccd1 vccd1 _14380_/C sky130_fd_sc_hd__clkinv_4
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08782_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08821_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07733_ _15333_/Q _15315_/Q vssd1 vssd1 vccd1 vccd1 _07734_/B sky130_fd_sc_hd__xor2_4
XFILLER_38_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07664_ _15205_/Q _07658_/C _14095_/B vssd1 vssd1 vccd1 vccd1 _07665_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09403_ _15366_/Q _09577_/B _09403_/C vssd1 vssd1 vccd1 vccd1 _09414_/A sky130_fd_sc_hd__and3_1
XFILLER_80_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09334_ _15355_/Q _09334_/B _09334_/C vssd1 vssd1 vccd1 vccd1 _09334_/Y sky130_fd_sc_hd__nand3_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09265_ _09266_/B _09266_/C _09266_/A vssd1 vssd1 vccd1 vccd1 _09267_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08216_ _08217_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08218_/A sky130_fd_sc_hd__nor2_1
X_09196_ _09196_/A vssd1 vssd1 vccd1 vccd1 _09211_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08147_ _08147_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _08264_/A sky130_fd_sc_hd__xnor2_4
XFILLER_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08078_ _12763_/A _07799_/B _08077_/X vssd1 vssd1 vccd1 vccd1 _08222_/B sky130_fd_sc_hd__o21a_1
XFILLER_134_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10040_ _10047_/A _10038_/Y _10039_/Y _10035_/C vssd1 vssd1 vccd1 vccd1 _10042_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11991_ _15770_/Q _12107_/B _12000_/C vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__and3_1
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ _13730_/A _13730_/B _13734_/A vssd1 vssd1 vccd1 vccd1 _16054_/D sky130_fd_sc_hd__nor3_1
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10942_ _10939_/X _10941_/Y _10936_/B _10937_/C vssd1 vssd1 vccd1 vccd1 _10944_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_83_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ _13659_/A _13659_/B _13660_/X vssd1 vssd1 vccd1 vccd1 _16041_/D sky130_fd_sc_hd__a21oi_1
X_10873_ _11507_/A vssd1 vssd1 vccd1 vccd1 _11161_/B sky130_fd_sc_hd__buf_2
XFILLER_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15400_ _15483_/CLK _15400_/D vssd1 vssd1 vccd1 vccd1 _15400_/Q sky130_fd_sc_hd__dfxtp_1
X_12612_ _12610_/Y _12605_/C _12607_/X _12608_/Y vssd1 vssd1 vccd1 vccd1 _12613_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13592_ _16031_/Q _13794_/B _13597_/C vssd1 vssd1 vccd1 vccd1 _13592_/Y sky130_fd_sc_hd__nand3_1
X_15331_ _15339_/CLK _15331_/D vssd1 vssd1 vccd1 vccd1 _15331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12543_ _12543_/A _12543_/B _12543_/C vssd1 vssd1 vccd1 vccd1 _12544_/C sky130_fd_sc_hd__nand3_1
XFILLER_40_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15262_ _15282_/CLK _15262_/D vssd1 vssd1 vccd1 vccd1 _15262_/Q sky130_fd_sc_hd__dfxtp_2
X_12474_ _12510_/A _12474_/B _12474_/C vssd1 vssd1 vccd1 vccd1 _12475_/A sky130_fd_sc_hd__and3_1
X_14213_ _14343_/A _14213_/B _14213_/C vssd1 vssd1 vccd1 vccd1 _14214_/A sky130_fd_sc_hd__and3_1
X_16372__21 vssd1 vssd1 vccd1 vccd1 _16372__21/HI io_oeb[4] sky130_fd_sc_hd__conb_1
X_11425_ _12569_/A vssd1 vssd1 vccd1 vccd1 _11425_/X sky130_fd_sc_hd__clkbuf_2
X_15193_ _07710_/X _15191_/A _15192_/Y vssd1 vssd1 vccd1 vccd1 _16367_/D sky130_fd_sc_hd__o21a_1
XANTENNA_7 _12758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14144_ _14364_/A vssd1 vssd1 vccd1 vccd1 _14320_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11356_ _11353_/X _11354_/Y _11355_/Y _11351_/C vssd1 vssd1 vccd1 vccd1 _11358_/B
+ sky130_fd_sc_hd__o211ai_1
X_10307_ _10301_/B _10302_/C _10304_/X _10305_/Y vssd1 vssd1 vccd1 vccd1 _10308_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14075_ _16120_/Q _14080_/C _07634_/A vssd1 vssd1 vccd1 vccd1 _14077_/C sky130_fd_sc_hd__a21o_1
X_11287_ _11309_/A _11287_/B _11287_/C vssd1 vssd1 vccd1 vccd1 _11288_/A sky130_fd_sc_hd__and3_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _13026_/A _13026_/B vssd1 vssd1 vccd1 vccd1 _13031_/C sky130_fd_sc_hd__nor2_1
X_10238_ _15496_/Q _10276_/C _10181_/X vssd1 vssd1 vccd1 vccd1 _10240_/B sky130_fd_sc_hd__a21oi_1
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10169_ _10169_/A vssd1 vssd1 vccd1 vccd1 _10404_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14977_ _16319_/Q _14977_/B _14981_/C vssd1 vssd1 vccd1 vccd1 _14984_/A sky130_fd_sc_hd__and3_1
XFILLER_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13928_ _14328_/A vssd1 vssd1 vccd1 vccd1 _14413_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13859_ _13857_/A _13857_/B _13858_/X vssd1 vssd1 vccd1 vccd1 _16077_/D sky130_fd_sc_hd__a21oi_1
XFILLER_23_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15529_ _15655_/CLK _15529_/D vssd1 vssd1 vccd1 vccd1 _15529_/Q sky130_fd_sc_hd__dfxtp_1
X_09050_ _09058_/A _09050_/B _09050_/C vssd1 vssd1 vccd1 vccd1 _09051_/A sky130_fd_sc_hd__and3_1
XFILLER_129_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08001_ _08187_/A _08187_/B vssd1 vssd1 vccd1 vccd1 _08188_/A sky130_fd_sc_hd__xnor2_2
XFILLER_128_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09952_ _15452_/Q _10010_/B _09958_/C vssd1 vssd1 vccd1 vccd1 _09955_/B sky130_fd_sc_hd__nand3_1
X_08903_ _15279_/Q vssd1 vssd1 vccd1 vccd1 _08919_/C sky130_fd_sc_hd__clkinv_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09997_/A _09883_/B _09883_/C vssd1 vssd1 vccd1 vccd1 _09886_/B sky130_fd_sc_hd__or3_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08834_/A _08834_/B vssd1 vssd1 vccd1 vccd1 _08835_/B sky130_fd_sc_hd__nor2_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08765_ _08765_/A _08765_/B _08765_/C vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__and3_1
X_07716_ _15234_/Q vssd1 vssd1 vccd1 vccd1 _08610_/C sky130_fd_sc_hd__inv_2
XFILLER_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08696_ _08694_/Y _08690_/C _08692_/X _08693_/Y vssd1 vssd1 vccd1 vccd1 _08697_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_53_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07647_ _13275_/A vssd1 vssd1 vccd1 vccd1 _10950_/C sky130_fd_sc_hd__buf_4
XFILLER_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09317_ _15353_/Q _09354_/C _09316_/X vssd1 vssd1 vccd1 vccd1 _09319_/B sky130_fd_sc_hd__a21oi_1
X_09248_ _09472_/A _09251_/C vssd1 vssd1 vccd1 vccd1 _09248_/X sky130_fd_sc_hd__or2_1
X_09179_ _15332_/Q _09354_/B _09179_/C vssd1 vssd1 vccd1 vccd1 _09190_/B sky130_fd_sc_hd__and3_1
XFILLER_135_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11210_ _11249_/A _11210_/B _11210_/C vssd1 vssd1 vccd1 vccd1 _11211_/A sky130_fd_sc_hd__and3_1
X_12190_ _12226_/A _12190_/B _12190_/C vssd1 vssd1 vccd1 vccd1 _12191_/A sky130_fd_sc_hd__and3_1
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11141_ _11139_/Y _11133_/C _11146_/A _11138_/Y vssd1 vssd1 vccd1 vccd1 _11146_/B
+ sky130_fd_sc_hd__a211oi_1
X_11072_ _15626_/Q _11078_/C _10897_/X vssd1 vssd1 vccd1 vccd1 _11072_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_122_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10023_ _15463_/Q _10024_/C _09794_/X vssd1 vssd1 vccd1 vccd1 _10023_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14900_ _14905_/C vssd1 vssd1 vccd1 vccd1 _14916_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15880_ _15907_/CLK _15880_/D vssd1 vssd1 vccd1 vccd1 _15880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14831_ _14831_/A vssd1 vssd1 vccd1 vccd1 _16280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14762_ _14757_/A _14760_/B _14646_/X vssd1 vssd1 vccd1 vccd1 _14769_/C sky130_fd_sc_hd__o21a_1
XFILLER_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11974_ _11975_/B _11975_/C _11975_/A vssd1 vssd1 vccd1 vccd1 _11976_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13713_ _13713_/A _13716_/C vssd1 vssd1 vccd1 vccd1 _13713_/X sky130_fd_sc_hd__or2_1
X_10925_ _15602_/Q vssd1 vssd1 vccd1 vccd1 _10939_/B sky130_fd_sc_hd__inv_2
X_14693_ _14853_/A _14811_/B _14693_/C vssd1 vssd1 vccd1 vccd1 _14697_/A sky130_fd_sc_hd__and3_1
XFILLER_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13644_ _13641_/X _13642_/Y _13643_/Y _13638_/C vssd1 vssd1 vccd1 vccd1 _13646_/B
+ sky130_fd_sc_hd__o211ai_1
X_10856_ _15592_/Q _10855_/C _10624_/X vssd1 vssd1 vccd1 vccd1 _10857_/B sky130_fd_sc_hd__a21oi_1
XFILLER_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16364_/CLK _16363_/D vssd1 vssd1 vccd1 vccd1 _16363_/Q sky130_fd_sc_hd__dfxtp_2
X_13575_ _16029_/Q _13675_/B _13575_/C vssd1 vssd1 vccd1 vccd1 _13580_/A sky130_fd_sc_hd__and3_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10783_/X _10784_/Y _10786_/Y _10781_/C vssd1 vssd1 vccd1 vccd1 _10789_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15314_ _15356_/CLK _15314_/D vssd1 vssd1 vccd1 vccd1 _15314_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12526_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12565_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16294_ _16321_/CLK _16294_/D vssd1 vssd1 vccd1 vccd1 _16294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15245_ _15254_/CLK _15245_/D vssd1 vssd1 vccd1 vccd1 _15245_/Q sky130_fd_sc_hd__dfxtp_1
X_12457_ _15843_/Q _12462_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12457_/Y sky130_fd_sc_hd__a21oi_1
X_11408_ _15679_/Q _11409_/C _11237_/X vssd1 vssd1 vccd1 vccd1 _11408_/Y sky130_fd_sc_hd__a21oi_1
X_15176_ _16367_/Q _15176_/B _15176_/C vssd1 vssd1 vccd1 vccd1 _15178_/A sky130_fd_sc_hd__and3_1
XFILLER_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12388_ _12386_/Y _12381_/C _12383_/X _12385_/Y vssd1 vssd1 vccd1 vccd1 _12389_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ _14132_/A _14126_/Y _14122_/B _14123_/C vssd1 vssd1 vccd1 vccd1 _14129_/B
+ sky130_fd_sc_hd__o211a_1
X_11339_ _11373_/A _11339_/B _11343_/A vssd1 vssd1 vccd1 vccd1 _15666_/D sky130_fd_sc_hd__nor3_1
XFILLER_98_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ _14325_/A vssd1 vssd1 vccd1 vccd1 _14058_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13009_ _15932_/Q _13064_/B _13016_/C vssd1 vssd1 vccd1 vccd1 _13009_/X sky130_fd_sc_hd__and3_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08550_ _15236_/Q _08588_/C _07623_/X vssd1 vssd1 vccd1 vccd1 _08553_/B sky130_fd_sc_hd__a21oi_1
XFILLER_63_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08481_ hold3/X _13474_/A _08493_/C vssd1 vssd1 vccd1 vccd1 _08488_/A sky130_fd_sc_hd__and3_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09102_ _15320_/Q _09158_/B _09105_/C vssd1 vssd1 vccd1 vccd1 _09102_/X sky130_fd_sc_hd__and3_1
XFILLER_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09033_ _15309_/Q _09146_/B _09039_/C vssd1 vssd1 vccd1 vccd1 _09036_/B sky130_fd_sc_hd__nand3_1
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09935_ _09935_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09939_/C sky130_fd_sc_hd__nor2_1
XFILLER_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09866_ _09866_/A vssd1 vssd1 vccd1 vccd1 _15436_/D sky130_fd_sc_hd__clkbuf_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08817_ _15276_/Q _08823_/C _08575_/X vssd1 vssd1 vccd1 vccd1 _08817_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09797_ _09793_/X _09795_/Y _09796_/Y _09790_/C vssd1 vssd1 vccd1 vccd1 _09799_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08748_ _08742_/B _08743_/C _08745_/X _08746_/Y vssd1 vssd1 vccd1 vccd1 _08749_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _15255_/Q _08853_/B _08686_/C vssd1 vssd1 vccd1 vccd1 _08682_/B sky130_fd_sc_hd__nand3_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10710_/A _10710_/B _10710_/C vssd1 vssd1 vccd1 vccd1 _10711_/C sky130_fd_sc_hd__nand3_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _15723_/Q _11697_/C _11519_/X vssd1 vssd1 vccd1 vccd1 _11690_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ _10665_/C vssd1 vssd1 vccd1 vccd1 _10679_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13360_ _13410_/A _13360_/B _13360_/C vssd1 vssd1 vccd1 vccd1 _13361_/A sky130_fd_sc_hd__and3_1
X_10572_ _10572_/A _10572_/B vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__nor2_1
X_12311_ _15821_/Q _12369_/B _12317_/C vssd1 vssd1 vccd1 vccd1 _12314_/B sky130_fd_sc_hd__nand3_1
XFILLER_127_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13291_ _15979_/Q _13394_/B _13291_/C vssd1 vssd1 vccd1 vccd1 _13300_/A sky130_fd_sc_hd__and3_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15030_ _15030_/A vssd1 vssd1 vccd1 vccd1 _15106_/A sky130_fd_sc_hd__clkbuf_2
X_12242_ _12413_/A vssd1 vssd1 vccd1 vccd1 _12281_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _15798_/Q _12178_/C _12001_/X vssd1 vssd1 vccd1 vccd1 _12173_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11124_ _11133_/A _11124_/B _11124_/C vssd1 vssd1 vccd1 vccd1 _11125_/A sky130_fd_sc_hd__and3_1
XFILLER_96_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11055_ _11076_/A _11055_/B _11055_/C vssd1 vssd1 vccd1 vccd1 _11056_/A sky130_fd_sc_hd__and3_1
X_15932_ _15196_/Q _15932_/D vssd1 vssd1 vccd1 vccd1 _15932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _15460_/Q _10043_/C _09893_/X vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__a21oi_1
XFILLER_37_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15863_ _15961_/CLK _15863_/D vssd1 vssd1 vccd1 vccd1 _15863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14814_ _14814_/A vssd1 vssd1 vccd1 vccd1 _14814_/X sky130_fd_sc_hd__clkbuf_2
X_15794_ _15794_/CLK _15794_/D vssd1 vssd1 vccd1 vccd1 _15794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14745_ _16266_/Q _14743_/C _14744_/X vssd1 vssd1 vccd1 vccd1 _14747_/C sky130_fd_sc_hd__a21o_1
X_11957_ _12129_/A vssd1 vssd1 vccd1 vccd1 _11997_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10908_ _10906_/Y _10902_/C _10914_/A _10905_/Y vssd1 vssd1 vccd1 vccd1 _10914_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_60_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14676_ _14716_/A _14676_/B _14680_/B vssd1 vssd1 vccd1 vccd1 _16245_/D sky130_fd_sc_hd__nor3_1
X_11888_ _11894_/A _11886_/Y _11887_/Y _11883_/C vssd1 vssd1 vccd1 vccd1 _11890_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13627_ _13730_/A _13627_/B _13631_/A vssd1 vssd1 vccd1 vccd1 _16036_/D sky130_fd_sc_hd__nor3_1
XFILLER_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10839_ _10839_/A vssd1 vssd1 vccd1 vccd1 _15588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16346_ _16352_/CLK _16346_/D vssd1 vssd1 vccd1 vccd1 _16346_/Q sky130_fd_sc_hd__dfxtp_1
X_13558_ _13558_/A _13558_/B vssd1 vssd1 vccd1 vccd1 _13561_/C sky130_fd_sc_hd__nor2_1
XFILLER_146_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12509_ _12507_/Y _12503_/C _12505_/X _12506_/Y vssd1 vssd1 vccd1 vccd1 _12510_/C
+ sky130_fd_sc_hd__a211o_1
X_16277_ _16321_/CLK _16277_/D vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
X_13489_ _13489_/A vssd1 vssd1 vccd1 vccd1 _16011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15228_ _15230_/CLK _15228_/D vssd1 vssd1 vccd1 vccd1 _15228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15159_ _15013_/X _15157_/A _15158_/Y vssd1 vssd1 vccd1 vccd1 _16358_/D sky130_fd_sc_hd__o21a_1
XFILLER_141_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07981_ _10002_/A _07924_/B _07980_/X vssd1 vssd1 vccd1 vccd1 _08180_/B sky130_fd_sc_hd__o21a_1
XFILLER_99_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09720_ _09775_/A _09720_/B _09724_/A vssd1 vssd1 vccd1 vccd1 _15414_/D sky130_fd_sc_hd__nor3_1
XFILLER_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09651_ _09825_/A vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08602_ _08648_/A _08602_/B _08602_/C vssd1 vssd1 vccd1 vccd1 _08603_/A sky130_fd_sc_hd__and3_1
X_09582_ _09588_/A _09578_/Y _09581_/Y _09575_/C vssd1 vssd1 vccd1 vccd1 _09584_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08533_ _15233_/Q _08532_/C _13715_/A vssd1 vssd1 vccd1 vccd1 _08534_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08464_ _08465_/A _08465_/C _08465_/B vssd1 vssd1 vccd1 vccd1 _08466_/B sky130_fd_sc_hd__o21ai_1
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08395_ _15212_/Q vssd1 vssd1 vccd1 vccd1 _08397_/A sky130_fd_sc_hd__inv_2
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09016_ _10169_/A vssd1 vssd1 vccd1 vccd1 _09250_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09918_ _10785_/A vssd1 vssd1 vccd1 vccd1 _10150_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09849_ _09847_/X _09848_/Y _09843_/B _09844_/C vssd1 vssd1 vccd1 vccd1 _09851_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12860_ _12934_/A _12860_/B _12864_/B vssd1 vssd1 vccd1 vccd1 _15905_/D sky130_fd_sc_hd__nor3_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _15742_/Q _11811_/B _11814_/C vssd1 vssd1 vccd1 vccd1 _11811_/X sky130_fd_sc_hd__and3_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _15896_/Q _12954_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__and3_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14524_/Y _14527_/X _14529_/Y vssd1 vssd1 vccd1 vccd1 _16211_/D sky130_fd_sc_hd__o21a_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11742_/A _11742_/B _11742_/C vssd1 vssd1 vccd1 vccd1 _11743_/C sky130_fd_sc_hd__nand3_1
XFILLER_54_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14461_/A _14461_/B vssd1 vssd1 vccd1 vccd1 _16196_/D sky130_fd_sc_hd__nor2_1
X_11673_ _11673_/A vssd1 vssd1 vccd1 vccd1 _15718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16200_ _16247_/CLK _16200_/D vssd1 vssd1 vccd1 vccd1 _16200_/Q sky130_fd_sc_hd__dfxtp_2
X_13412_ _13666_/A vssd1 vssd1 vccd1 vccd1 _13412_/X sky130_fd_sc_hd__clkbuf_2
X_10624_ _11488_/A vssd1 vssd1 vccd1 vccd1 _10624_/X sky130_fd_sc_hd__clkbuf_4
X_14392_ _14386_/B _14387_/C _14397_/A _14390_/Y vssd1 vssd1 vccd1 vccd1 _14397_/B
+ sky130_fd_sc_hd__a211oi_1
X_16131_ _16142_/CLK _16131_/D vssd1 vssd1 vccd1 vccd1 _16131_/Q sky130_fd_sc_hd__dfxtp_1
X_13343_ _15988_/Q _13349_/C _13342_/X vssd1 vssd1 vccd1 vccd1 _13343_/Y sky130_fd_sc_hd__a21oi_1
X_10555_ _15545_/Q _10561_/C _10318_/X vssd1 vssd1 vccd1 vccd1 _10555_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16062_ _16129_/CLK _16062_/D vssd1 vssd1 vccd1 vccd1 _16062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ _13274_/A vssd1 vssd1 vccd1 vccd1 _15974_/D sky130_fd_sc_hd__clkbuf_1
X_10486_ _10484_/X _10485_/Y _10481_/B _10482_/C vssd1 vssd1 vccd1 vccd1 _10488_/B
+ sky130_fd_sc_hd__o211ai_1
X_15013_ _15013_/A vssd1 vssd1 vccd1 vccd1 _15013_/X sky130_fd_sc_hd__buf_2
XFILLER_136_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12225_ _12223_/Y _12219_/C _12221_/X _12222_/Y vssd1 vssd1 vccd1 vccd1 _12226_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_123_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12156_ _12726_/A vssd1 vssd1 vccd1 vccd1 _12383_/B sky130_fd_sc_hd__clkbuf_2
X_11107_ _15632_/Q _11221_/B _11113_/C vssd1 vssd1 vccd1 vccd1 _11110_/B sky130_fd_sc_hd__nand3_1
X_12087_ _15785_/Q _12092_/C _12086_/X vssd1 vssd1 vccd1 vccd1 _12089_/C sky130_fd_sc_hd__a21o_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11038_ _12188_/A vssd1 vssd1 vccd1 vccd1 _11038_/X sky130_fd_sc_hd__clkbuf_2
X_15915_ _07603_/A _15915_/D vssd1 vssd1 vccd1 vccd1 _15915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15846_ _15907_/CLK _15846_/D vssd1 vssd1 vccd1 vccd1 _15846_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15777_ _15794_/CLK _15777_/D vssd1 vssd1 vccd1 vccd1 _15777_/Q sky130_fd_sc_hd__dfxtp_1
X_12989_ _13077_/A _12989_/B _12993_/A vssd1 vssd1 vccd1 vccd1 _15927_/D sky130_fd_sc_hd__nor3_1
XFILLER_17_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14728_ _14765_/A _14731_/C vssd1 vssd1 vccd1 vccd1 _14730_/A sky130_fd_sc_hd__and2_1
XFILLER_60_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14659_ _16259_/Q _16258_/Q hold9/X _14620_/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__o31a_4
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08180_ _08180_/A _08180_/B vssd1 vssd1 vccd1 vccd1 _08180_/Y sky130_fd_sc_hd__nor2_1
X_16329_ _16337_/CLK _16329_/D vssd1 vssd1 vccd1 vccd1 _16329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07964_ _08198_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07975_/A sky130_fd_sc_hd__nor2_4
X_09703_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09704_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07895_ _15324_/Q vssd1 vssd1 vccd1 vccd1 _09196_/A sky130_fd_sc_hd__inv_2
XFILLER_110_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09634_ _09632_/Y _09626_/C _09628_/X _09629_/Y vssd1 vssd1 vccd1 vccd1 _09635_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09565_ _15390_/Q _09623_/B _09565_/C vssd1 vssd1 vccd1 vccd1 _09565_/Y sky130_fd_sc_hd__nand3_1
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08516_ _15230_/Q _10957_/C _08522_/C vssd1 vssd1 vccd1 vccd1 _08516_/Y sky130_fd_sc_hd__nand3_1
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09496_ _15381_/Q _09496_/B _09496_/C vssd1 vssd1 vccd1 vccd1 _09496_/X sky130_fd_sc_hd__and3_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08447_ _08446_/A _08446_/B _14363_/A vssd1 vssd1 vccd1 vccd1 _08448_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ _08378_/A _08378_/B vssd1 vssd1 vccd1 vccd1 _08379_/A sky130_fd_sc_hd__and2_1
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ _10404_/A vssd1 vssd1 vccd1 vccd1 _10386_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10271_ _15500_/Q _10391_/B _10276_/C vssd1 vssd1 vccd1 vccd1 _10271_/Y sky130_fd_sc_hd__nand3_1
XFILLER_105_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _12010_/A _12010_/B vssd1 vssd1 vccd1 vccd1 _12011_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13961_ _13956_/Y _13959_/X _13960_/Y vssd1 vssd1 vccd1 vccd1 _16094_/D sky130_fd_sc_hd__o21a_1
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15700_ _15763_/CLK _15700_/D vssd1 vssd1 vccd1 vccd1 _15700_/Q sky130_fd_sc_hd__dfxtp_1
X_12912_ _12910_/Y _12906_/C _12917_/A _12909_/Y vssd1 vssd1 vccd1 vccd1 _12917_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13892_ _14261_/A vssd1 vssd1 vccd1 vccd1 _14598_/B sky130_fd_sc_hd__buf_2
X_15631_ _15194_/Q _15631_/D vssd1 vssd1 vccd1 vccd1 _15631_/Q sky130_fd_sc_hd__dfxtp_1
X_12843_ _12851_/A _12843_/B _12843_/C vssd1 vssd1 vccd1 vccd1 _12844_/A sky130_fd_sc_hd__and3_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ _15655_/CLK _15562_/D vssd1 vssd1 vccd1 vccd1 _15562_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12774_/A _12774_/B _12774_/C vssd1 vssd1 vccd1 vccd1 _12775_/C sky130_fd_sc_hd__nand3_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _16212_/Q _14593_/B _14513_/C vssd1 vssd1 vccd1 vccd1 _14520_/A sky130_fd_sc_hd__and3_1
X_11725_ _11723_/A _11723_/B _11724_/X vssd1 vssd1 vccd1 vccd1 _15726_/D sky130_fd_sc_hd__a21oi_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _15224_/Q _15493_/D vssd1 vssd1 vccd1 vccd1 _15493_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14444_ _14443_/X _14442_/Y _14309_/X vssd1 vssd1 vccd1 vccd1 _14444_/Y sky130_fd_sc_hd__a21oi_1
X_11656_ _15717_/Q _11662_/C _11425_/X vssd1 vssd1 vccd1 vccd1 _11656_/Y sky130_fd_sc_hd__a21oi_1
X_10607_ _10615_/A _10607_/B _10607_/C vssd1 vssd1 vccd1 vccd1 _10608_/A sky130_fd_sc_hd__and3_1
X_14375_ _16196_/Q _16195_/Q _16194_/Q _14202_/X vssd1 vssd1 vccd1 vccd1 _16179_/D
+ sky130_fd_sc_hd__o31a_1
X_11587_ _11585_/Y _11580_/C _11583_/X _11584_/Y vssd1 vssd1 vccd1 vccd1 _11588_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16114_ _16114_/CLK _16114_/D vssd1 vssd1 vccd1 vccd1 _16114_/Q sky130_fd_sc_hd__dfxtp_1
X_13326_ _13326_/A vssd1 vssd1 vccd1 vccd1 _15983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ _10559_/A _10538_/B _10538_/C vssd1 vssd1 vccd1 vccd1 _10539_/A sky130_fd_sc_hd__and3_1
X_16045_ _16050_/CLK _16045_/D vssd1 vssd1 vccd1 vccd1 _16045_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ _13281_/A _13257_/B _13257_/C vssd1 vssd1 vccd1 vccd1 _13258_/A sky130_fd_sc_hd__and3_1
X_10469_ _15530_/Q vssd1 vssd1 vccd1 vccd1 _10484_/C sky130_fd_sc_hd__inv_2
XFILLER_142_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12208_ _15804_/Q _12434_/B _12208_/C vssd1 vssd1 vccd1 vccd1 _12208_/X sky130_fd_sc_hd__and3_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13188_ _15961_/Q _13193_/C _14605_/B vssd1 vssd1 vccd1 vccd1 _13188_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12139_ _12172_/C vssd1 vssd1 vccd1 vccd1 _12178_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07680_ input6/X vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15829_ _07603_/A _15829_/D vssd1 vssd1 vccd1 vccd1 _15829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09350_ _15357_/Q _09524_/B _09354_/C vssd1 vssd1 vccd1 vccd1 _09350_/Y sky130_fd_sc_hd__nand3_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08301_ _08301_/A _08301_/B vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09281_ _09288_/A _09281_/B _09281_/C vssd1 vssd1 vccd1 vccd1 _09282_/A sky130_fd_sc_hd__and3_1
X_08232_ _08301_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08233_/B sky130_fd_sc_hd__or2_2
XFILLER_21_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08163_ _08163_/A _08163_/B vssd1 vssd1 vccd1 vccd1 _08429_/C sky130_fd_sc_hd__xor2_4
XFILLER_119_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08094_ _10289_/A _10177_/A _08093_/Y vssd1 vssd1 vccd1 vccd1 _08096_/B sky130_fd_sc_hd__o21a_1
XFILLER_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08996_ _15302_/Q _08996_/B _09001_/C vssd1 vssd1 vccd1 vccd1 _08996_/Y sky130_fd_sc_hd__nand3_1
XFILLER_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07947_ _07633_/C _07929_/B _07928_/B vssd1 vssd1 vccd1 vccd1 _08159_/A sky130_fd_sc_hd__o21ai_4
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07878_ _16017_/Q _16035_/Q vssd1 vssd1 vccd1 vccd1 _07879_/B sky130_fd_sc_hd__or2_1
X_09617_ _09615_/X _09616_/Y _09612_/B _09613_/C vssd1 vssd1 vccd1 vccd1 _09619_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_71_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09548_ _15388_/Q _09663_/B _09557_/C vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__and3_1
XFILLER_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09479_ _09479_/A vssd1 vssd1 vccd1 vccd1 _15376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _15695_/Q _11510_/B _11518_/C vssd1 vssd1 vccd1 vccd1 _11515_/B sky130_fd_sc_hd__nand3_1
X_12490_ _12490_/A vssd1 vssd1 vccd1 vccd1 _15847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11441_ _11477_/A _11441_/B _11441_/C vssd1 vssd1 vccd1 vccd1 _11442_/A sky130_fd_sc_hd__and3_1
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ _14379_/A vssd1 vssd1 vccd1 vccd1 _14337_/B sky130_fd_sc_hd__buf_2
X_11372_ _11370_/Y _11365_/C _11377_/A _11368_/Y vssd1 vssd1 vccd1 vccd1 _11377_/B
+ sky130_fd_sc_hd__a211oi_1
X_13111_ _15950_/Q _13109_/C _14869_/A vssd1 vssd1 vccd1 vccd1 _13111_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_125_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10323_ _10323_/A _10323_/B _10323_/C vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__and3_1
X_14091_ _14123_/A _14091_/B _14091_/C vssd1 vssd1 vccd1 vccd1 _14092_/A sky130_fd_sc_hd__and3_1
XFILLER_106_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13042_ _15938_/Q _13078_/C _13041_/X vssd1 vssd1 vccd1 vccd1 _13044_/B sky130_fd_sc_hd__a21oi_1
X_10254_ _15499_/Q _10256_/C _10083_/X vssd1 vssd1 vccd1 vccd1 _10254_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10185_ _15488_/Q _10298_/B _10191_/C vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__nand3_1
XFILLER_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14993_ _14993_/A vssd1 vssd1 vccd1 vccd1 _15142_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13944_ _13944_/A vssd1 vssd1 vccd1 vccd1 _16091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13875_ _13980_/A _13875_/B _13881_/A vssd1 vssd1 vccd1 vccd1 _16081_/D sky130_fd_sc_hd__nor3_1
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15614_ _15194_/Q _15614_/D vssd1 vssd1 vccd1 vccd1 _15614_/Q sky130_fd_sc_hd__dfxtp_1
X_12826_ _15902_/Q _12935_/B _12832_/C vssd1 vssd1 vccd1 vccd1 _12829_/B sky130_fd_sc_hd__nand3_1
X_15545_ _15655_/CLK _15545_/D vssd1 vssd1 vccd1 vccd1 _15545_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12869_/A _12757_/B _12757_/C vssd1 vssd1 vccd1 vccd1 _12760_/B sky130_fd_sc_hd__or3_1
XFILLER_91_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11708_/A _11708_/B _11708_/C vssd1 vssd1 vccd1 vccd1 _11709_/A sky130_fd_sc_hd__and3_1
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15476_ _15485_/CLK _15476_/D vssd1 vssd1 vccd1 vccd1 _15476_/Q sky130_fd_sc_hd__dfxtp_1
X_12688_ _12686_/Y _12680_/C _12693_/A _12685_/Y vssd1 vssd1 vccd1 vccd1 _12693_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14427_ _14427_/A _14427_/B _14431_/A vssd1 vssd1 vccd1 vccd1 _16189_/D sky130_fd_sc_hd__nor3_1
X_11639_ _11653_/A _11639_/B _11639_/C vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__and3_1
X_14358_ _16178_/Q _14357_/C _14270_/X vssd1 vssd1 vccd1 vccd1 _14359_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13309_ _13154_/X _13307_/C _13206_/X vssd1 vssd1 vccd1 vccd1 _13309_/Y sky130_fd_sc_hd__o21ai_1
X_14289_ _16165_/Q _14337_/B _14289_/C vssd1 vssd1 vccd1 vccd1 _14295_/A sky130_fd_sc_hd__and3_1
XFILLER_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16028_ _16031_/CLK _16028_/D vssd1 vssd1 vccd1 vccd1 _16028_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_143_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08850_ _10007_/A vssd1 vssd1 vccd1 vccd1 _09088_/B sky130_fd_sc_hd__clkbuf_2
X_07801_ _16152_/Q vssd1 vssd1 vccd1 vccd1 _14289_/C sky130_fd_sc_hd__inv_2
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08781_ _08779_/A _08779_/B _08780_/X vssd1 vssd1 vccd1 vccd1 _15268_/D sky130_fd_sc_hd__a21oi_1
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07732_ _16332_/Q vssd1 vssd1 vccd1 vccd1 _08109_/A sky130_fd_sc_hd__inv_2
XFILLER_84_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07663_ _15176_/B vssd1 vssd1 vccd1 vccd1 _14095_/B sky130_fd_sc_hd__buf_4
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09402_ _09402_/A vssd1 vssd1 vccd1 vccd1 _15364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09333_ _15356_/Q _09334_/C _09220_/X vssd1 vssd1 vccd1 vccd1 _09333_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09264_ _15345_/Q _09270_/C _09205_/X vssd1 vssd1 vccd1 vccd1 _09266_/C sky130_fd_sc_hd__a21o_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ _08037_/A _08037_/B _08214_/X vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__a21oi_1
X_09195_ _15350_/Q _15349_/Q _15348_/Q _09194_/X vssd1 vssd1 vccd1 vccd1 _15333_/D
+ sky130_fd_sc_hd__o31a_1
X_08146_ _08260_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__xor2_4
XFILLER_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08077_ _12874_/A _08077_/B vssd1 vssd1 vccd1 vccd1 _08077_/X sky130_fd_sc_hd__or2_1
XFILLER_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_08979_ _11229_/A vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__buf_4
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11990_ _11990_/A vssd1 vssd1 vccd1 vccd1 _15768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10941_ _15606_/Q _10950_/B _10940_/X vssd1 vssd1 vccd1 vccd1 _10941_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13660_ _13713_/A _13662_/C vssd1 vssd1 vccd1 vccd1 _13660_/X sky130_fd_sc_hd__or2_1
XFILLER_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10872_ _15595_/Q _10910_/C _10760_/X vssd1 vssd1 vccd1 vccd1 _10875_/B sky130_fd_sc_hd__a21oi_1
X_12611_ _12607_/X _12608_/Y _12610_/Y _12605_/C vssd1 vssd1 vccd1 vccd1 _12613_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13591_ _14300_/A vssd1 vssd1 vccd1 vccd1 _13794_/B sky130_fd_sc_hd__buf_2
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15330_ _15337_/CLK _15330_/D vssd1 vssd1 vccd1 vccd1 _15330_/Q sky130_fd_sc_hd__dfxtp_1
X_12542_ _12543_/B _12543_/C _12543_/A vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ _15359_/CLK _15261_/D vssd1 vssd1 vccd1 vccd1 _15261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12473_ _12471_/B _12471_/C _12472_/X vssd1 vssd1 vccd1 vccd1 _12474_/C sky130_fd_sc_hd__o21ai_1
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14212_ _14212_/A _14212_/B _14212_/C vssd1 vssd1 vccd1 vccd1 _14213_/C sky130_fd_sc_hd__nand3_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11424_ _11424_/A vssd1 vssd1 vccd1 vccd1 _12569_/A sky130_fd_sc_hd__clkbuf_4
X_15192_ _13926_/X _15191_/A _14054_/A vssd1 vssd1 vccd1 vccd1 _15192_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_8 _14466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14363_/A vssd1 vssd1 vccd1 vccd1 _14321_/A sky130_fd_sc_hd__clkbuf_2
X_11355_ _15669_/Q _11409_/B _11355_/C vssd1 vssd1 vccd1 vccd1 _11355_/Y sky130_fd_sc_hd__nand3_1
XFILLER_99_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _10304_/X _10305_/Y _10301_/B _10302_/C vssd1 vssd1 vccd1 vccd1 _10308_/B
+ sky130_fd_sc_hd__o211ai_1
X_14074_ _16120_/Q _14074_/B _14080_/C vssd1 vssd1 vccd1 vccd1 _14077_/B sky130_fd_sc_hd__nand3_1
X_11286_ _11286_/A _11286_/B _11286_/C vssd1 vssd1 vccd1 vccd1 _11287_/C sky130_fd_sc_hd__nand3_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13025_ _13025_/A _13025_/B vssd1 vssd1 vccd1 vccd1 _13026_/B sky130_fd_sc_hd__nor2_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _10268_/C vssd1 vssd1 vccd1 vccd1 _10276_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_67_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10168_ _10166_/A _10166_/B _10167_/X vssd1 vssd1 vccd1 vccd1 _15483_/D sky130_fd_sc_hd__a21oi_1
X_10099_ _10388_/A vssd1 vssd1 vccd1 vccd1 _10219_/A sky130_fd_sc_hd__buf_2
X_14976_ _16319_/Q _14994_/C _14901_/X vssd1 vssd1 vccd1 vccd1 _14978_/B sky130_fd_sc_hd__a21oi_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13927_ _13925_/X _13917_/B _13926_/X vssd1 vssd1 vccd1 vccd1 _13932_/A sky130_fd_sc_hd__a21oi_1
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _14644_/A _13861_/C vssd1 vssd1 vccd1 vccd1 _13858_/X sky130_fd_sc_hd__or2_1
XFILLER_90_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12809_ _12809_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _12813_/C sky130_fd_sc_hd__nor2_1
X_13789_ _13789_/A _13789_/B _13789_/C vssd1 vssd1 vccd1 vccd1 _13790_/A sky130_fd_sc_hd__and3_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15528_ _15655_/CLK _15528_/D vssd1 vssd1 vccd1 vccd1 _15528_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15459_ _15483_/CLK _15459_/D vssd1 vssd1 vccd1 vccd1 _15459_/Q sky130_fd_sc_hd__dfxtp_2
X_08000_ _08209_/A _08000_/B vssd1 vssd1 vccd1 vccd1 _08187_/B sky130_fd_sc_hd__and2_1
XFILLER_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09951_ _10064_/A _09951_/B _09955_/A vssd1 vssd1 vccd1 vccd1 _15450_/D sky130_fd_sc_hd__nor3_1
XFILLER_131_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08902_ hold29/X _15304_/Q _15303_/Q _08901_/X vssd1 vssd1 vccd1 vccd1 _15288_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _10114_/A vssd1 vssd1 vccd1 vccd1 _09922_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _08839_/B _08833_/B vssd1 vssd1 vccd1 vccd1 _08835_/A sky130_fd_sc_hd__or2_1
XFILLER_112_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08762_/Y _08756_/C _08758_/X _08759_/Y vssd1 vssd1 vccd1 vccd1 _08765_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07715_ _15207_/Q vssd1 vssd1 vccd1 vccd1 _07945_/A sky130_fd_sc_hd__inv_2
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08695_ _08692_/X _08693_/Y _08694_/Y _08690_/C vssd1 vssd1 vccd1 vccd1 _08697_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07646_ _12661_/A vssd1 vssd1 vccd1 vccd1 _13275_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09316_ _10181_/A vssd1 vssd1 vccd1 vccd1 _09316_/X sky130_fd_sc_hd__buf_2
XFILLER_22_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09247_ _09247_/A _09247_/B vssd1 vssd1 vccd1 vccd1 _09251_/C sky130_fd_sc_hd__nor2_1
XFILLER_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09178_ _09202_/A _09178_/B _09183_/B vssd1 vssd1 vccd1 vccd1 _15330_/D sky130_fd_sc_hd__nor3_1
X_08129_ _07729_/A _07729_/B _08128_/X vssd1 vssd1 vccd1 vccd1 _08244_/B sky130_fd_sc_hd__o21a_1
X_11140_ _11146_/A _11138_/Y _11139_/Y _11133_/C vssd1 vssd1 vccd1 vccd1 _11142_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11071_ _15626_/Q _11244_/B _11078_/C vssd1 vssd1 vccd1 vccd1 _11071_/X sky130_fd_sc_hd__and3_1
XFILLER_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10022_ _15463_/Q _10022_/B _10024_/C vssd1 vssd1 vccd1 vccd1 _10022_/X sky130_fd_sc_hd__and3_1
XFILLER_76_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14830_ _14946_/A _14830_/B _14830_/C vssd1 vssd1 vccd1 vccd1 _14831_/A sky130_fd_sc_hd__and3_1
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11973_ _15767_/Q _11978_/C _11798_/X vssd1 vssd1 vccd1 vccd1 _11975_/C sky130_fd_sc_hd__a21o_1
X_14761_ _14759_/A _14759_/B _14760_/X vssd1 vssd1 vccd1 vccd1 _16264_/D sky130_fd_sc_hd__a21oi_1
XFILLER_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10924_ _15610_/Q _15609_/Q _15608_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _15602_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_72_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13712_ _13712_/A _13712_/B vssd1 vssd1 vccd1 vccd1 _13716_/C sky130_fd_sc_hd__nor2_1
XFILLER_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14692_ _15005_/A vssd1 vssd1 vccd1 vccd1 _14853_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13643_ _16040_/Q _13794_/B _13648_/C vssd1 vssd1 vccd1 vccd1 _13643_/Y sky130_fd_sc_hd__nand3_1
X_10855_ _15592_/Q _11143_/B _10855_/C vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__and3_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13574_ _16029_/Q _13605_/C _13573_/X vssd1 vssd1 vccd1 vccd1 _13576_/B sky130_fd_sc_hd__a21oi_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _16362_/CLK _16362_/D vssd1 vssd1 vccd1 vccd1 _16362_/Q sky130_fd_sc_hd__dfxtp_2
X_10786_ _15580_/Q _11073_/B _10792_/C vssd1 vssd1 vccd1 vccd1 _10786_/Y sky130_fd_sc_hd__nand3_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _15322_/CLK _15313_/D vssd1 vssd1 vccd1 vccd1 _15313_/Q sky130_fd_sc_hd__dfxtp_1
X_12525_ _12523_/A _12523_/B _12524_/X vssd1 vssd1 vccd1 vccd1 _15852_/D sky130_fd_sc_hd__a21oi_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16293_ _16321_/CLK _16293_/D vssd1 vssd1 vccd1 vccd1 _16293_/Q sky130_fd_sc_hd__dfxtp_1
X_15244_ _15254_/CLK _15244_/D vssd1 vssd1 vccd1 vccd1 _15244_/Q sky130_fd_sc_hd__dfxtp_2
X_12456_ _15843_/Q _12512_/B _12456_/C vssd1 vssd1 vccd1 vccd1 _12465_/A sky130_fd_sc_hd__and3_1
XFILLER_126_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11407_ _15679_/Q _11525_/B _11409_/C vssd1 vssd1 vccd1 vccd1 _11407_/X sky130_fd_sc_hd__and3_1
X_15175_ _15175_/A _15175_/B _15179_/B vssd1 vssd1 vccd1 vccd1 _16362_/D sky130_fd_sc_hd__nor3_1
X_12387_ _12383_/X _12385_/Y _12386_/Y _12381_/C vssd1 vssd1 vccd1 vccd1 _12389_/B
+ sky130_fd_sc_hd__o211ai_1
X_14126_ _16131_/Q _14125_/C _14033_/X vssd1 vssd1 vccd1 vccd1 _14126_/Y sky130_fd_sc_hd__a21oi_1
X_11338_ _15667_/Q _11449_/B _11347_/C vssd1 vssd1 vccd1 vccd1 _11343_/A sky130_fd_sc_hd__and3_1
XFILLER_99_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14057_ _13920_/X _14054_/B _14056_/Y vssd1 vssd1 vccd1 vccd1 _16114_/D sky130_fd_sc_hd__o21a_1
X_11269_ _11268_/B _11268_/C _11038_/X vssd1 vssd1 vccd1 vccd1 _11270_/C sky130_fd_sc_hd__o21ai_1
XFILLER_97_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13008_ _13008_/A vssd1 vssd1 vccd1 vccd1 _15930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14959_ _14957_/A _14957_/B _14958_/X vssd1 vssd1 vccd1 vccd1 _16309_/D sky130_fd_sc_hd__a21oi_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08480_ _12650_/A vssd1 vssd1 vccd1 vccd1 _13474_/A sky130_fd_sc_hd__buf_6
XFILLER_35_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09101_ _09101_/A vssd1 vssd1 vccd1 vccd1 _15318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09032_ _09066_/A _09032_/B _09036_/A vssd1 vssd1 vccd1 vccd1 _15307_/D sky130_fd_sc_hd__nor3_1
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _09934_/A _09934_/B vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09865_ _09865_/A _09865_/B _09865_/C vssd1 vssd1 vccd1 vccd1 _09866_/A sky130_fd_sc_hd__and3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _15276_/Q _08872_/B _08823_/C vssd1 vssd1 vccd1 vccd1 _08816_/X sky130_fd_sc_hd__and3_1
X_09796_ _15426_/Q _09911_/B _09796_/C vssd1 vssd1 vccd1 vccd1 _09796_/Y sky130_fd_sc_hd__nand3_1
XFILLER_39_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08747_ _08745_/X _08746_/Y _08742_/B _08743_/C vssd1 vssd1 vccd1 vccd1 _08749_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08774_/A _08678_/B _08682_/A vssd1 vssd1 vccd1 vccd1 _15253_/D sky130_fd_sc_hd__nor3_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07629_ _10354_/A vssd1 vssd1 vccd1 vccd1 _13045_/B sky130_fd_sc_hd__buf_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10654_/C vssd1 vssd1 vccd1 vccd1 _10665_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10571_ _10577_/B _10571_/B vssd1 vssd1 vccd1 vccd1 _10573_/A sky130_fd_sc_hd__or2_1
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ _12368_/A _12310_/B _12314_/A vssd1 vssd1 vccd1 vccd1 _15819_/D sky130_fd_sc_hd__nor3_1
X_13290_ _13290_/A vssd1 vssd1 vccd1 vccd1 _15976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12241_ _12239_/A _12239_/B _12240_/X vssd1 vssd1 vccd1 vccd1 _15807_/D sky130_fd_sc_hd__a21oi_1
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ _15798_/Q _12228_/B _12172_/C vssd1 vssd1 vccd1 vccd1 _12181_/A sky130_fd_sc_hd__and3_1
XFILLER_122_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11123_ _11121_/Y _11117_/C _11119_/X _11120_/Y vssd1 vssd1 vccd1 vccd1 _11124_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_123_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11054_ _11054_/A _11054_/B _11054_/C vssd1 vssd1 vccd1 vccd1 _11055_/C sky130_fd_sc_hd__nand3_1
XFILLER_77_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15931_ _15196_/Q _15931_/D vssd1 vssd1 vccd1 vccd1 _15931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10005_ _10037_/C vssd1 vssd1 vccd1 vccd1 _10043_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15862_ _15907_/CLK _15862_/D vssd1 vssd1 vccd1 vccd1 _15862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14813_ _14813_/A _14813_/B vssd1 vssd1 vccd1 vccd1 _16276_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15793_ _15794_/CLK _15793_/D vssd1 vssd1 vccd1 vccd1 _15793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14744_ _14980_/A vssd1 vssd1 vccd1 vccd1 _14744_/X sky130_fd_sc_hd__clkbuf_2
X_11956_ _11954_/A _11954_/B _11955_/X vssd1 vssd1 vccd1 vccd1 _15762_/D sky130_fd_sc_hd__a21oi_1
XFILLER_83_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10907_ _10914_/A _10905_/Y _10906_/Y _10902_/C vssd1 vssd1 vccd1 vccd1 _10909_/B
+ sky130_fd_sc_hd__o211a_1
X_11887_ _15752_/Q _11887_/B _11891_/C vssd1 vssd1 vccd1 vccd1 _11887_/Y sky130_fd_sc_hd__nand3_1
X_14675_ _14668_/B _14669_/C _14680_/A _14673_/Y vssd1 vssd1 vccd1 vccd1 _14680_/B
+ sky130_fd_sc_hd__a211oi_1
X_13626_ _16038_/Q _13675_/B _13626_/C vssd1 vssd1 vccd1 vccd1 _13631_/A sky130_fd_sc_hd__and3_1
X_10838_ _10845_/A _10838_/B _10838_/C vssd1 vssd1 vccd1 vccd1 _10839_/A sky130_fd_sc_hd__and3_1
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ _16358_/CLK _16345_/D vssd1 vssd1 vccd1 vccd1 _16345_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10769_ _10769_/A vssd1 vssd1 vccd1 vccd1 _15577_/D sky130_fd_sc_hd__clkbuf_1
X_13557_ _13557_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13558_/B sky130_fd_sc_hd__nor2_1
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12508_ _12505_/X _12506_/Y _12507_/Y _12503_/C vssd1 vssd1 vccd1 vccd1 _12510_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_146_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16276_ _16321_/CLK _16276_/D vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfxtp_1
X_13488_ _13538_/A _13488_/B _13488_/C vssd1 vssd1 vccd1 vccd1 _13489_/A sky130_fd_sc_hd__and3_1
XFILLER_145_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15227_ _15230_/CLK _15227_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
X_12439_ _12439_/A vssd1 vssd1 vccd1 vccd1 _15839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15158_ _13926_/X _15157_/A _15014_/X vssd1 vssd1 vccd1 vccd1 _15158_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14109_ _14109_/A vssd1 vssd1 vccd1 vccd1 _16123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07980_ _10121_/A _07980_/B vssd1 vssd1 vccd1 vccd1 _07980_/X sky130_fd_sc_hd__or2_1
X_15089_ _14970_/X _15088_/A _15014_/X vssd1 vssd1 vccd1 vccd1 _15089_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ _09648_/A _09648_/B _09649_/X vssd1 vssd1 vccd1 vccd1 _15402_/D sky130_fd_sc_hd__a21oi_1
X_08601_ _08600_/B _08600_/C _08541_/X vssd1 vssd1 vccd1 vccd1 _08602_/C sky130_fd_sc_hd__o21ai_1
XFILLER_94_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09581_ _15392_/Q _09813_/B _09585_/C vssd1 vssd1 vccd1 vccd1 _09581_/Y sky130_fd_sc_hd__nand3_1
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08532_ _15233_/Q _08775_/B _08532_/C vssd1 vssd1 vccd1 vccd1 _08540_/B sky130_fd_sc_hd__and3_1
XFILLER_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08463_ _08468_/A _08468_/B vssd1 vssd1 vccd1 vccd1 _08465_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08394_ _15212_/Q _08403_/B _08452_/B vssd1 vssd1 vccd1 vccd1 _08411_/A sky130_fd_sc_hd__a21oi_2
Xclkbuf_leaf_30_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _16100_/CLK sky130_fd_sc_hd__clkbuf_16
X_09015_ _14163_/A vssd1 vssd1 vccd1 vccd1 _10169_/A sky130_fd_sc_hd__buf_4
XFILLER_128_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09917_ _15446_/Q _09925_/C _09741_/X vssd1 vssd1 vccd1 vccd1 _09917_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_97_clk _15665_/CLK vssd1 vssd1 vccd1 vccd1 _15701_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09848_ _15435_/Q _09855_/C _09786_/X vssd1 vssd1 vccd1 vccd1 _09848_/Y sky130_fd_sc_hd__a21oi_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ _15425_/Q _09784_/C _09778_/X vssd1 vssd1 vccd1 vccd1 _09781_/C sky130_fd_sc_hd__a21o_1
XFILLER_74_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11810_/A vssd1 vssd1 vccd1 vccd1 _15740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12790_/A vssd1 vssd1 vccd1 vccd1 _15894_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11741_ _11742_/B _11742_/C _11742_/A vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__a21o_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11672_ _11708_/A _11672_/B _11672_/C vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__and3_1
XFILLER_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14328_/X _14372_/X _14454_/B _14459_/X vssd1 vssd1 vccd1 vccd1 _14461_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _15556_/Q _10798_/B _10623_/C vssd1 vssd1 vccd1 vccd1 _10634_/B sky130_fd_sc_hd__and3_1
X_13411_ _13411_/A vssd1 vssd1 vccd1 vccd1 _15997_/D sky130_fd_sc_hd__clkbuf_1
X_14391_ _14397_/A _14390_/Y _14386_/B _14387_/C vssd1 vssd1 vccd1 vccd1 _14393_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _16060_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16130_ _16142_/CLK _16130_/D vssd1 vssd1 vccd1 vccd1 _16130_/Q sky130_fd_sc_hd__dfxtp_1
X_13342_ _13598_/A vssd1 vssd1 vccd1 vccd1 _13342_/X sky130_fd_sc_hd__buf_2
X_10554_ _15545_/Q _10609_/B _10561_/C vssd1 vssd1 vccd1 vccd1 _10554_/X sky130_fd_sc_hd__and3_1
XFILLER_6_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13273_ _13281_/A _13273_/B _13273_/C vssd1 vssd1 vccd1 vccd1 _13274_/A sky130_fd_sc_hd__and3_1
XFILLER_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16061_ _16124_/CLK _16061_/D vssd1 vssd1 vccd1 vccd1 _16061_/Q sky130_fd_sc_hd__dfxtp_1
X_10485_ _15534_/Q _10492_/C _10364_/X vssd1 vssd1 vccd1 vccd1 _10485_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12224_ _12221_/X _12222_/Y _12223_/Y _12219_/C vssd1 vssd1 vccd1 vccd1 _12226_/B
+ sky130_fd_sc_hd__o211ai_1
X_15012_ _15012_/A _15012_/B vssd1 vssd1 vccd1 vccd1 _16321_/D sky130_fd_sc_hd__nor2_1
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12155_ _12155_/A vssd1 vssd1 vccd1 vccd1 _15794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11106_ _11220_/A _11106_/B _11110_/A vssd1 vssd1 vccd1 vccd1 _15630_/D sky130_fd_sc_hd__nor3_1
XFILLER_110_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12086_ _12654_/A vssd1 vssd1 vccd1 vccd1 _12086_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_88_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15351_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11037_ _11037_/A vssd1 vssd1 vccd1 vccd1 _12188_/A sky130_fd_sc_hd__clkbuf_4
X_15914_ _15196_/Q _15914_/D vssd1 vssd1 vccd1 vccd1 _15914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15845_ _15845_/CLK _15845_/D vssd1 vssd1 vccd1 vccd1 _15845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15776_ _15794_/CLK _15776_/D vssd1 vssd1 vccd1 vccd1 _15776_/Q sky130_fd_sc_hd__dfxtp_1
X_12988_ _15928_/Q _13043_/B _12996_/C vssd1 vssd1 vccd1 vccd1 _12993_/A sky130_fd_sc_hd__and3_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14727_ _07675_/X _14720_/A _14723_/B _14726_/Y vssd1 vssd1 vccd1 vccd1 _16256_/D
+ sky130_fd_sc_hd__o31a_1
X_11939_ _11936_/X _11937_/Y _11938_/Y _11934_/C vssd1 vssd1 vccd1 vccd1 _11941_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14658_ _07707_/X _14656_/A _14657_/Y vssd1 vssd1 vccd1 vccd1 _16241_/D sky130_fd_sc_hd__o21a_1
XFILLER_60_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _13609_/A _13609_/B vssd1 vssd1 vccd1 vccd1 _13613_/C sky130_fd_sc_hd__nor2_1
X_14589_ _14590_/B _14590_/C _14590_/A vssd1 vssd1 vccd1 vccd1 _14591_/B sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_12_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _16007_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16328_ _16344_/CLK _16328_/D vssd1 vssd1 vccd1 vccd1 _16328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16259_ _16268_/CLK _16259_/D vssd1 vssd1 vccd1 vccd1 _16259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07963_ _07963_/A _07963_/B _07963_/C vssd1 vssd1 vccd1 vccd1 _07964_/B sky130_fd_sc_hd__and3_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_79_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15377_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09702_ _09708_/B _09702_/B vssd1 vssd1 vccd1 vccd1 _09704_/A sky130_fd_sc_hd__or2_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07894_ _15306_/Q _08152_/B vssd1 vssd1 vccd1 vccd1 _07935_/A sky130_fd_sc_hd__xnor2_4
XFILLER_68_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09633_ _09628_/X _09629_/Y _09632_/Y _09626_/C vssd1 vssd1 vccd1 vccd1 _09635_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09564_ _15391_/Q _09565_/C _09506_/X vssd1 vssd1 vccd1 vccd1 _09564_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08515_ _12847_/A vssd1 vssd1 vccd1 vccd1 _10957_/C sky130_fd_sc_hd__buf_2
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _09495_/A vssd1 vssd1 vccd1 vccd1 _15379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08446_ _08446_/A _08446_/B vssd1 vssd1 vccd1 vccd1 _08448_/A sky130_fd_sc_hd__or2_1
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08377_ _08375_/A _08375_/B _14363_/A vssd1 vssd1 vccd1 vccd1 _08378_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10270_ _15501_/Q _10276_/C _10269_/X vssd1 vssd1 vccd1 vccd1 _10270_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13960_ _13956_/Y _13959_/X _13922_/X vssd1 vssd1 vccd1 vccd1 _13960_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _12917_/A _12909_/Y _12910_/Y _12906_/C vssd1 vssd1 vccd1 vccd1 _12913_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13891_ _16087_/Q _13950_/B _13903_/C vssd1 vssd1 vccd1 vccd1 _13896_/A sky130_fd_sc_hd__and3_1
XFILLER_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15630_ _15194_/Q _15630_/D vssd1 vssd1 vccd1 vccd1 _15630_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _12840_/Y _12836_/C _12838_/X _12839_/Y vssd1 vssd1 vccd1 vccd1 _12843_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15655_/CLK _15561_/D vssd1 vssd1 vccd1 vccd1 _15561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12774_/B _12774_/C _12774_/A vssd1 vssd1 vccd1 vccd1 _12775_/B sky130_fd_sc_hd__a21o_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14512_/A vssd1 vssd1 vccd1 vccd1 _16208_/D sky130_fd_sc_hd__clkbuf_1
X_11724_ _11780_/A _11727_/C vssd1 vssd1 vccd1 vccd1 _11724_/X sky130_fd_sc_hd__or2_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _15224_/Q _15492_/D vssd1 vssd1 vccd1 vccd1 _15492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _15717_/Q _11655_/B _11655_/C vssd1 vssd1 vccd1 vccd1 _11665_/A sky130_fd_sc_hd__and3_1
X_14443_ _14443_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14443_/X sky130_fd_sc_hd__or2_1
X_10606_ _10604_/Y _10600_/C _10602_/X _10603_/Y vssd1 vssd1 vccd1 vccd1 _10607_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11586_ _11583_/X _11584_/Y _11585_/Y _11580_/C vssd1 vssd1 vccd1 vccd1 _11588_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_128_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14374_ _14374_/A _14374_/B vssd1 vssd1 vccd1 vccd1 _16178_/D sky130_fd_sc_hd__nor2_1
X_16113_ _16114_/CLK _16113_/D vssd1 vssd1 vccd1 vccd1 _16113_/Q sky130_fd_sc_hd__dfxtp_1
X_10537_ _10537_/A _10537_/B _10537_/C vssd1 vssd1 vccd1 vccd1 _10538_/C sky130_fd_sc_hd__nand3_1
X_13325_ _13339_/A _13325_/B _13325_/C vssd1 vssd1 vccd1 vccd1 _13326_/A sky130_fd_sc_hd__and3_1
XFILLER_127_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _16124_/CLK _16044_/D vssd1 vssd1 vccd1 vccd1 _16044_/Q sky130_fd_sc_hd__dfxtp_1
X_10468_ _15538_/Q _15537_/Q _15536_/Q _10409_/X vssd1 vssd1 vccd1 vccd1 _15530_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_89_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13256_ _13255_/B _13255_/C _14892_/A vssd1 vssd1 vccd1 vccd1 _13257_/C sky130_fd_sc_hd__o21ai_1
XFILLER_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12207_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12434_/B sky130_fd_sc_hd__clkbuf_2
X_13187_ _15961_/Q _13394_/B _13187_/C vssd1 vssd1 vccd1 vccd1 _13197_/A sky130_fd_sc_hd__and3_1
X_10399_ _13250_/A vssd1 vssd1 vccd1 vccd1 _11551_/A sky130_fd_sc_hd__buf_2
XFILLER_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12138_ _12159_/C vssd1 vssd1 vccd1 vccd1 _12172_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12069_ _12067_/A _12067_/B _12068_/X vssd1 vssd1 vccd1 vccd1 _15780_/D sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_1_clk _15665_/CLK vssd1 vssd1 vccd1 vccd1 _15890_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15828_ _07603_/A _15828_/D vssd1 vssd1 vccd1 vccd1 _15828_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15759_ _15794_/CLK _15759_/D vssd1 vssd1 vccd1 vccd1 _15759_/Q sky130_fd_sc_hd__dfxtp_1
X_08300_ _08233_/B _08300_/B vssd1 vssd1 vccd1 vccd1 _08301_/B sky130_fd_sc_hd__and2b_1
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09280_ _09278_/Y _09274_/C _09276_/X _09277_/Y vssd1 vssd1 vccd1 vccd1 _09281_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08231_ _08231_/A _08231_/B _08231_/C vssd1 vssd1 vccd1 vccd1 _08232_/B sky130_fd_sc_hd__and3_1
XFILLER_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08162_ _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08163_/B sky130_fd_sc_hd__xor2_4
XFILLER_119_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08093_ _15521_/Q _08093_/B vssd1 vssd1 vccd1 vccd1 _08093_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08995_ _15303_/Q _09001_/C _08873_/X vssd1 vssd1 vccd1 vccd1 _08995_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07946_ _08421_/A _07946_/B _07946_/C vssd1 vssd1 vccd1 vccd1 _15206_/D sky130_fd_sc_hd__nor3_1
XFILLER_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ _16017_/Q _16035_/Q vssd1 vssd1 vccd1 vccd1 _07879_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09616_ _15399_/Q _09623_/C _09497_/X vssd1 vssd1 vccd1 vccd1 _09616_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09547_ _15388_/Q _09585_/C _09316_/X vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__a21oi_1
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _09519_/A _09478_/B _09478_/C vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__and3_1
XFILLER_52_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08429_ state1[2] _08433_/A _08429_/C vssd1 vssd1 vccd1 vccd1 _08429_/X sky130_fd_sc_hd__and3_1
XFILLER_8_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11440_ _11439_/B _11439_/C _11327_/X vssd1 vssd1 vccd1 vccd1 _11441_/C sky130_fd_sc_hd__o21ai_1
XFILLER_50_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11371_ _11377_/A _11368_/Y _11370_/Y _11365_/C vssd1 vssd1 vccd1 vccd1 _11373_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10322_ _10320_/Y _10315_/C _10317_/X _10319_/Y vssd1 vssd1 vccd1 vccd1 _10323_/C
+ sky130_fd_sc_hd__a211o_1
X_13110_ _13534_/A vssd1 vssd1 vccd1 vccd1 _14869_/A sky130_fd_sc_hd__clkbuf_4
X_14090_ _14088_/Y _14084_/C _14086_/X _14087_/Y vssd1 vssd1 vccd1 vccd1 _14091_/C
+ sky130_fd_sc_hd__a211o_1
X_13041_ _13041_/A vssd1 vssd1 vccd1 vccd1 _13041_/X sky130_fd_sc_hd__clkbuf_4
X_10253_ _15499_/Q _10310_/B _10256_/C vssd1 vssd1 vccd1 vccd1 _10253_/X sky130_fd_sc_hd__and3_1
XFILLER_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10184_ _10219_/A _10184_/B _10188_/A vssd1 vssd1 vccd1 vccd1 _15486_/D sky130_fd_sc_hd__nor3_1
XFILLER_132_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14992_ _15023_/A hold31/X _14997_/B vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__nor3_1
X_13943_ _14029_/A _13943_/B _13943_/C vssd1 vssd1 vccd1 vccd1 _13944_/A sky130_fd_sc_hd__and3_1
XFILLER_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13874_ _16084_/Q _14117_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13881_/A sky130_fd_sc_hd__and3_1
XFILLER_47_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15613_ _15194_/Q _15613_/D vssd1 vssd1 vccd1 vccd1 _15613_/Q sky130_fd_sc_hd__dfxtp_1
X_12825_ _12934_/A _12825_/B _12829_/A vssd1 vssd1 vccd1 vccd1 _15900_/D sky130_fd_sc_hd__nor3_1
X_15544_ _15655_/CLK _15544_/D vssd1 vssd1 vccd1 vccd1 _15544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12796_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11705_/Y _11700_/C _11702_/X _11703_/Y vssd1 vssd1 vccd1 vccd1 _11708_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _15484_/CLK _15475_/D vssd1 vssd1 vccd1 vccd1 _15475_/Q sky130_fd_sc_hd__dfxtp_1
X_12687_ _12693_/A _12685_/Y _12686_/Y _12680_/C vssd1 vssd1 vccd1 vccd1 _12689_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14426_ _16192_/Q _14546_/B _14426_/C vssd1 vssd1 vccd1 vccd1 _14431_/A sky130_fd_sc_hd__and3_1
X_11638_ _11631_/B _11632_/C _11635_/X _11636_/Y vssd1 vssd1 vccd1 vccd1 _11639_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14357_ _16178_/Q _14357_/B _14357_/C vssd1 vssd1 vccd1 vccd1 _14357_/X sky130_fd_sc_hd__and3_1
XFILLER_128_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11569_ _11569_/A vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13308_ _13308_/A vssd1 vssd1 vccd1 vccd1 _15979_/D sky130_fd_sc_hd__clkbuf_1
X_14288_ _16165_/Q _14313_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14290_/B sky130_fd_sc_hd__a21oi_1
X_16027_ _16040_/CLK _16027_/D vssd1 vssd1 vccd1 vccd1 _16027_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13239_ _13239_/A vssd1 vssd1 vccd1 vccd1 _13348_/A sky130_fd_sc_hd__buf_2
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07800_ _11388_/A _07800_/B vssd1 vssd1 vccd1 vccd1 _08044_/A sky130_fd_sc_hd__xnor2_1
X_08780_ _08893_/A _08783_/C vssd1 vssd1 vccd1 vccd1 _08780_/X sky130_fd_sc_hd__or2_1
XFILLER_85_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07731_ _16314_/Q vssd1 vssd1 vccd1 vccd1 _07737_/A sky130_fd_sc_hd__inv_2
X_07662_ _13130_/A vssd1 vssd1 vccd1 vccd1 _15176_/B sky130_fd_sc_hd__buf_4
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09401_ _09401_/A _09401_/B _09401_/C vssd1 vssd1 vccd1 vccd1 _09402_/A sky130_fd_sc_hd__and3_1
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09332_ _15356_/Q _09444_/B _09334_/C vssd1 vssd1 vccd1 vccd1 _09332_/X sky130_fd_sc_hd__and3_1
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09263_ _15345_/Q _09432_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09266_/B sky130_fd_sc_hd__nand3_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08214_ _08036_/B _08214_/B vssd1 vssd1 vccd1 vccd1 _08214_/X sky130_fd_sc_hd__and2b_1
X_09194_ _09541_/A vssd1 vssd1 vccd1 vccd1 _09194_/X sky130_fd_sc_hd__buf_4
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08145_ _07828_/A _07828_/B _08144_/Y vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__o21a_1
XFILLER_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08076_ _08227_/B _08305_/B vssd1 vssd1 vccd1 vccd1 _08222_/A sky130_fd_sc_hd__xor2_1
XFILLER_146_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08978_ _08978_/A vssd1 vssd1 vccd1 vccd1 _15299_/D sky130_fd_sc_hd__clkbuf_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07929_ _07929_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _07930_/B sky130_fd_sc_hd__xnor2_4
XFILLER_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10940_ _10940_/A vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ _10904_/C vssd1 vssd1 vccd1 vccd1 _10910_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12610_ _15867_/Q _12840_/B _12610_/C vssd1 vssd1 vccd1 vccd1 _12610_/Y sky130_fd_sc_hd__nand3_1
X_13590_ _16032_/Q _13597_/C _13437_/X vssd1 vssd1 vccd1 vccd1 _13590_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12541_ _15857_/Q _12546_/C _12370_/X vssd1 vssd1 vccd1 vccd1 _12543_/C sky130_fd_sc_hd__a21o_1
XFILLER_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15260_ _15260_/CLK _15260_/D vssd1 vssd1 vccd1 vccd1 _15260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12472_ _12758_/A vssd1 vssd1 vccd1 vccd1 _12472_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14211_ _14212_/B _14212_/C _14212_/A vssd1 vssd1 vccd1 vccd1 _14213_/B sky130_fd_sc_hd__a21o_1
X_11423_ _15681_/Q _11655_/B _11423_/C vssd1 vssd1 vccd1 vccd1 _11434_/A sky130_fd_sc_hd__and3_1
X_15191_ _15191_/A _15191_/B vssd1 vssd1 vccd1 vccd1 _16366_/D sky130_fd_sc_hd__nor2_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_9 _14466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _15670_/Q _11355_/C _11237_/X vssd1 vssd1 vccd1 vccd1 _11354_/Y sky130_fd_sc_hd__a21oi_1
X_14142_ _14136_/Y _14137_/X _14139_/B vssd1 vssd1 vccd1 vccd1 _14145_/B sky130_fd_sc_hd__o21a_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10305_ _15507_/Q _10312_/C _10075_/X vssd1 vssd1 vccd1 vccd1 _10305_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11285_ _11286_/B _11286_/C _11286_/A vssd1 vssd1 vccd1 vccd1 _11287_/B sky130_fd_sc_hd__a21o_1
X_14073_ _14073_/A vssd1 vssd1 vccd1 vccd1 _14123_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10236_ _10256_/C vssd1 vssd1 vccd1 vccd1 _10268_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13024_ _13031_/B _13024_/B vssd1 vssd1 vccd1 vccd1 _13026_/A sky130_fd_sc_hd__or2_1
XFILLER_140_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10167_ _10338_/A _10171_/C vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__or2_1
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10098_ _10098_/A vssd1 vssd1 vccd1 vccd1 _15472_/D sky130_fd_sc_hd__clkbuf_1
X_14975_ _14981_/C vssd1 vssd1 vccd1 vccd1 _14994_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13926_ _14326_/A vssd1 vssd1 vccd1 vccd1 _13926_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13857_ _13857_/A _13857_/B vssd1 vssd1 vccd1 vccd1 _13861_/C sky130_fd_sc_hd__nor2_1
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12808_ _12808_/A _12808_/B vssd1 vssd1 vccd1 vccd1 _12809_/B sky130_fd_sc_hd__nor2_1
X_13788_ _13782_/B _13783_/C _13785_/X _13786_/Y vssd1 vssd1 vccd1 vccd1 _13789_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15527_ _15655_/CLK _15527_/D vssd1 vssd1 vccd1 vccd1 _15527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _12737_/Y _12732_/C _12735_/X _12736_/Y vssd1 vssd1 vccd1 vccd1 _12740_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ _15485_/CLK _15458_/D vssd1 vssd1 vccd1 vccd1 _15458_/Q sky130_fd_sc_hd__dfxtp_1
X_14409_ _14401_/Y _14403_/X _14405_/B vssd1 vssd1 vccd1 vccd1 _14410_/B sky130_fd_sc_hd__o21a_1
X_15389_ _15484_/CLK _15389_/D vssd1 vssd1 vccd1 vccd1 _15389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09950_ _15451_/Q _09950_/B _09958_/C vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__and3_1
XFILLER_103_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08901_ _09541_/A vssd1 vssd1 vccd1 vccd1 _08901_/X sky130_fd_sc_hd__buf_2
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _10169_/A vssd1 vssd1 vccd1 vccd1 _10114_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08832_ _15278_/Q _08831_/C _08590_/X vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__a21oi_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08763_ _08758_/X _08759_/Y _08762_/Y _08756_/C vssd1 vssd1 vccd1 vccd1 _08765_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_73_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07714_ _07707_/X _07703_/A _07713_/Y vssd1 vssd1 vccd1 vccd1 _15205_/D sky130_fd_sc_hd__o21a_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08694_ _15256_/Q _08753_/B _08694_/C vssd1 vssd1 vccd1 vccd1 _08694_/Y sky130_fd_sc_hd__nand3_1
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07645_ _15204_/Q _14634_/B _07658_/C vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__and3_1
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09315_ _09348_/C vssd1 vssd1 vccd1 vccd1 _09354_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09246_ _10110_/A vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__clkbuf_2
X_09177_ _09175_/Y _09171_/C _09183_/A _09174_/Y vssd1 vssd1 vccd1 vccd1 _09183_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08128_ _15165_/C _08128_/B vssd1 vssd1 vccd1 vccd1 _08128_/X sky130_fd_sc_hd__or2_1
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08059_ _14466_/C _08059_/B vssd1 vssd1 vccd1 vccd1 _08059_/X sky130_fd_sc_hd__or2_1
XFILLER_122_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11070_ _11070_/A vssd1 vssd1 vccd1 vccd1 _15624_/D sky130_fd_sc_hd__clkbuf_1
X_10021_ _10021_/A vssd1 vssd1 vccd1 vccd1 _15461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14760_ _14843_/A _14760_/B vssd1 vssd1 vccd1 vccd1 _14760_/X sky130_fd_sc_hd__or2_1
X_11972_ _15767_/Q _12085_/B _11978_/C vssd1 vssd1 vccd1 vccd1 _11975_/B sky130_fd_sc_hd__nand3_1
X_13711_ _13711_/A _13711_/B vssd1 vssd1 vccd1 vccd1 _13712_/B sky130_fd_sc_hd__nor2_1
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10923_ _10923_/A vssd1 vssd1 vccd1 vccd1 _15601_/D sky130_fd_sc_hd__clkbuf_1
X_14691_ _14691_/A _14691_/B vssd1 vssd1 vccd1 vccd1 _16248_/D sky130_fd_sc_hd__nor2_1
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13642_ _16041_/Q _13648_/C _13437_/X vssd1 vssd1 vccd1 vccd1 _13642_/Y sky130_fd_sc_hd__a21oi_1
X_10854_ _11197_/A vssd1 vssd1 vccd1 vccd1 _11143_/B sky130_fd_sc_hd__buf_2
XFILLER_25_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16364_/CLK _16361_/D vssd1 vssd1 vccd1 vccd1 _16361_/Q sky130_fd_sc_hd__dfxtp_2
X_13573_ _14287_/A vssd1 vssd1 vccd1 vccd1 _13573_/X sky130_fd_sc_hd__buf_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _10785_/A vssd1 vssd1 vccd1 vccd1 _11073_/B sky130_fd_sc_hd__clkbuf_4
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15312_ _15312_/CLK _15312_/D vssd1 vssd1 vccd1 vccd1 _15312_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _12636_/A _12527_/C vssd1 vssd1 vccd1 vccd1 _12524_/X sky130_fd_sc_hd__or2_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _16304_/CLK _16292_/D vssd1 vssd1 vccd1 vccd1 _16292_/Q sky130_fd_sc_hd__dfxtp_1
X_15243_ _15260_/CLK _15243_/D vssd1 vssd1 vccd1 vccd1 _15243_/Q sky130_fd_sc_hd__dfxtp_2
X_12455_ _12455_/A vssd1 vssd1 vccd1 vccd1 _15841_/D sky130_fd_sc_hd__clkbuf_1
X_11406_ _11406_/A vssd1 vssd1 vccd1 vccd1 _15677_/D sky130_fd_sc_hd__clkbuf_1
X_15174_ _15168_/B _15169_/C _15179_/A _15172_/Y vssd1 vssd1 vccd1 vccd1 _15179_/B
+ sky130_fd_sc_hd__a211oi_1
X_12386_ _15831_/Q _12554_/B _12386_/C vssd1 vssd1 vccd1 vccd1 _12386_/Y sky130_fd_sc_hd__nand3_1
X_14125_ _16131_/Q _14256_/B _14125_/C vssd1 vssd1 vccd1 vccd1 _14132_/A sky130_fd_sc_hd__and3_1
X_11337_ _15667_/Q _11374_/C _11336_/X vssd1 vssd1 vccd1 vccd1 _11339_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14056_ _13921_/X _14054_/B _14049_/X vssd1 vssd1 vccd1 vccd1 _14056_/Y sky130_fd_sc_hd__a21oi_1
X_11268_ _11439_/A _11268_/B _11268_/C vssd1 vssd1 vccd1 vccd1 _11270_/B sky130_fd_sc_hd__or3_1
X_13007_ _13014_/A _13007_/B _13007_/C vssd1 vssd1 vccd1 vccd1 _13008_/A sky130_fd_sc_hd__and3_1
X_10219_ _10219_/A _10219_/B _10223_/B vssd1 vssd1 vccd1 vccd1 _15491_/D sky130_fd_sc_hd__nor3_1
XFILLER_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11199_ _11488_/A vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14958_ _15041_/A _14958_/B vssd1 vssd1 vccd1 vccd1 _14958_/X sky130_fd_sc_hd__or2_1
XFILLER_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13909_ _14364_/A vssd1 vssd1 vccd1 vccd1 _15005_/A sky130_fd_sc_hd__clkbuf_2
X_14889_ _14889_/A _14889_/B vssd1 vssd1 vccd1 vccd1 _16293_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09100_ _09115_/A _09100_/B _09100_/C vssd1 vssd1 vccd1 vccd1 _09101_/A sky130_fd_sc_hd__and3_1
XFILLER_149_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09031_ _15308_/Q _09088_/B _09039_/C vssd1 vssd1 vccd1 vccd1 _09036_/A sky130_fd_sc_hd__and3_1
XFILLER_148_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09933_ _09939_/B _09933_/B vssd1 vssd1 vccd1 vccd1 _09935_/A sky130_fd_sc_hd__or2_1
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09864_ _09862_/Y _09858_/C _09860_/X _09861_/Y vssd1 vssd1 vccd1 vccd1 _09865_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _08815_/A vssd1 vssd1 vccd1 vccd1 _15274_/D sky130_fd_sc_hd__clkbuf_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09795_ _15427_/Q _09796_/C _09794_/X vssd1 vssd1 vccd1 vccd1 _09795_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08746_ _15265_/Q _08753_/C _08625_/X vssd1 vssd1 vccd1 vccd1 _08746_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_73_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08677_ _15254_/Q _08794_/B _08686_/C vssd1 vssd1 vccd1 vccd1 _08682_/A sky130_fd_sc_hd__and3_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ input2/X vssd1 vssd1 vccd1 vccd1 _10354_/A sky130_fd_sc_hd__buf_4
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10570_ _15547_/Q _10569_/C _10333_/X vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ _15339_/Q _09236_/C _09166_/X vssd1 vssd1 vccd1 vccd1 _09229_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12240_ _12352_/A _12243_/C vssd1 vssd1 vccd1 vccd1 _12240_/X sky130_fd_sc_hd__or2_1
XFILLER_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12171_ _12171_/A vssd1 vssd1 vccd1 vccd1 _15796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11122_ _11119_/X _11120_/Y _11121_/Y _11117_/C vssd1 vssd1 vccd1 vccd1 _11124_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11053_ _11054_/B _11054_/C _11054_/A vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__a21o_1
X_15930_ _15196_/Q _15930_/D vssd1 vssd1 vccd1 vccd1 _15930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10004_ _10024_/C vssd1 vssd1 vccd1 vccd1 _10037_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15861_ _15907_/CLK _15861_/D vssd1 vssd1 vccd1 vccd1 _15861_/Q sky130_fd_sc_hd__dfxtp_1
X_14812_ _14694_/X _14810_/A _14808_/X vssd1 vssd1 vccd1 vccd1 _14813_/B sky130_fd_sc_hd__o21ai_1
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15792_ _15794_/CLK _15792_/D vssd1 vssd1 vccd1 vccd1 _15792_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14743_ _16266_/Q _14743_/B _14743_/C vssd1 vssd1 vccd1 vccd1 _14747_/B sky130_fd_sc_hd__nand3_1
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11955_ _12068_/A _11958_/C vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__or2_1
XFILLER_72_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10906_ _15599_/Q _11023_/B _10910_/C vssd1 vssd1 vccd1 vccd1 _10906_/Y sky130_fd_sc_hd__nand3_1
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _14680_/A _14673_/Y _14668_/B _14669_/C vssd1 vssd1 vccd1 vccd1 _14676_/B
+ sky130_fd_sc_hd__o211a_1
X_11886_ _15753_/Q _11891_/C _11713_/X vssd1 vssd1 vccd1 vccd1 _11886_/Y sky130_fd_sc_hd__a21oi_1
Xrepeater10 _07603_/A vssd1 vssd1 vccd1 vccd1 _15907_/CLK sky130_fd_sc_hd__buf_12
X_13625_ _16038_/Q _13655_/C _13573_/X vssd1 vssd1 vccd1 vccd1 _13627_/B sky130_fd_sc_hd__a21oi_1
X_10837_ _10835_/Y _10829_/C _10831_/X _10832_/Y vssd1 vssd1 vccd1 vccd1 _10838_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16344_ _16344_/CLK _16344_/D vssd1 vssd1 vccd1 vccd1 _16344_/Q sky130_fd_sc_hd__dfxtp_2
X_13556_ _13561_/B _13556_/B vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__or2_1
XFILLER_9_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10768_ _10789_/A _10768_/B _10768_/C vssd1 vssd1 vccd1 vccd1 _10769_/A sky130_fd_sc_hd__and3_1
XFILLER_118_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ _15850_/Q _12507_/B _12512_/C vssd1 vssd1 vccd1 vccd1 _12507_/Y sky130_fd_sc_hd__nand3_1
X_16275_ _16321_/CLK _16275_/D vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_1
X_13487_ _13480_/B _13481_/C _13484_/X _13485_/Y vssd1 vssd1 vccd1 vccd1 _13488_/C
+ sky130_fd_sc_hd__a211o_1
X_10699_ _15574_/Q _15573_/Q _15572_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _15566_/D
+ sky130_fd_sc_hd__o31a_1
X_15226_ _16242_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _15226_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12438_ _12454_/A _12438_/B _12438_/C vssd1 vssd1 vccd1 vccd1 _12439_/A sky130_fd_sc_hd__and3_1
X_15157_ _15157_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _16357_/D sky130_fd_sc_hd__nor2_1
XFILLER_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12369_ _15830_/Q _12369_/B _12376_/C vssd1 vssd1 vccd1 vccd1 _12373_/B sky130_fd_sc_hd__nand3_1
XFILLER_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ _14123_/A _14108_/B _14108_/C vssd1 vssd1 vccd1 vccd1 _14109_/A sky130_fd_sc_hd__and3_1
X_15088_ _15088_/A _15088_/B vssd1 vssd1 vccd1 vccd1 _16339_/D sky130_fd_sc_hd__nor2_1
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14039_ _16114_/Q _14046_/C _13893_/X vssd1 vssd1 vccd1 vccd1 _14041_/B sky130_fd_sc_hd__a21oi_1
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08600_ _08839_/A _08600_/B _08600_/C vssd1 vssd1 vccd1 vccd1 _08602_/B sky130_fd_sc_hd__or3_1
XFILLER_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09580_ _10736_/A vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__buf_2
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08531_ _09699_/A vssd1 vssd1 vccd1 vccd1 _08775_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08462_ state1[7] _08462_/B vssd1 vssd1 vccd1 vccd1 _08468_/B sky130_fd_sc_hd__and2_1
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ _08393_/A _08393_/B vssd1 vssd1 vccd1 vccd1 _08452_/B sky130_fd_sc_hd__xor2_4
XFILLER_149_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09014_ _09012_/A _09012_/B _09013_/X vssd1 vssd1 vccd1 vccd1 _15304_/D sky130_fd_sc_hd__a21oi_1
XFILLER_128_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09916_ _15446_/Q _10029_/B _09925_/C vssd1 vssd1 vccd1 vccd1 _09916_/X sky130_fd_sc_hd__and3_1
XFILLER_59_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09847_ _15435_/Q _10074_/B _09847_/C vssd1 vssd1 vccd1 vccd1 _09847_/X sky130_fd_sc_hd__and3_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09778_ _09778_/A vssd1 vssd1 vccd1 vccd1 _09778_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _08729_/A vssd1 vssd1 vccd1 vccd1 _15260_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _15731_/Q _11745_/C _11512_/X vssd1 vssd1 vccd1 vccd1 _11742_/C sky130_fd_sc_hd__a21o_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11670_/B _11670_/C _11615_/X vssd1 vssd1 vccd1 vccd1 _11672_/C sky130_fd_sc_hd__o21ai_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13410_/A _13410_/B _13410_/C vssd1 vssd1 vccd1 vccd1 _13411_/A sky130_fd_sc_hd__and3_1
X_10622_ _10645_/A _10622_/B _10627_/B vssd1 vssd1 vccd1 vccd1 _15554_/D sky130_fd_sc_hd__nor3_1
X_14390_ _16185_/Q _14389_/C _14300_/X vssd1 vssd1 vccd1 vccd1 _14390_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13341_ _15988_/Q _13394_/B _13341_/C vssd1 vssd1 vccd1 vccd1 _13352_/A sky130_fd_sc_hd__and3_1
X_10553_ _10553_/A vssd1 vssd1 vccd1 vccd1 _15543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16060_ _16060_/CLK _16060_/D vssd1 vssd1 vccd1 vccd1 _16060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13272_ _13272_/A _13272_/B _13272_/C vssd1 vssd1 vccd1 vccd1 _13273_/C sky130_fd_sc_hd__nand3_1
X_10484_ _15534_/Q _10654_/B _10484_/C vssd1 vssd1 vccd1 vccd1 _10484_/X sky130_fd_sc_hd__and3_1
XFILLER_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15011_ _14892_/X _15009_/A _15007_/X vssd1 vssd1 vccd1 vccd1 _15012_/B sky130_fd_sc_hd__o21ai_1
X_12223_ _15805_/Q _12223_/B _12228_/C vssd1 vssd1 vccd1 vccd1 _12223_/Y sky130_fd_sc_hd__nand3_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12154_ _12170_/A _12154_/B _12154_/C vssd1 vssd1 vccd1 vccd1 _12155_/A sky130_fd_sc_hd__and3_1
XFILLER_78_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11105_ _15631_/Q _11161_/B _11113_/C vssd1 vssd1 vccd1 vccd1 _11110_/A sky130_fd_sc_hd__and3_1
XFILLER_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12085_ _15785_/Q _12085_/B _12092_/C vssd1 vssd1 vccd1 vccd1 _12089_/B sky130_fd_sc_hd__nand3_1
XFILLER_78_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11036_ _11151_/A _11036_/B _11036_/C vssd1 vssd1 vccd1 vccd1 _11040_/B sky130_fd_sc_hd__or3_1
X_15913_ _07603_/A _15913_/D vssd1 vssd1 vccd1 vccd1 _15913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15844_ _15907_/CLK _15844_/D vssd1 vssd1 vccd1 vccd1 _15844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15775_ _15794_/CLK _15775_/D vssd1 vssd1 vccd1 vccd1 _15775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12987_ _15928_/Q _13022_/C _12767_/X vssd1 vssd1 vccd1 vccd1 _12989_/B sky130_fd_sc_hd__a21oi_1
XFILLER_92_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14726_ _14847_/A _14731_/C vssd1 vssd1 vccd1 vccd1 _14726_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11938_ _15760_/Q _11938_/B _11943_/C vssd1 vssd1 vccd1 vccd1 _11938_/Y sky130_fd_sc_hd__nand3_1
XFILLER_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14657_ _07710_/X _14656_/A _14614_/X vssd1 vssd1 vccd1 vccd1 _14657_/Y sky130_fd_sc_hd__a21oi_1
X_11869_ _12726_/A vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13608_ _13608_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13609_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14588_ _16229_/Q _14593_/C _07632_/A vssd1 vssd1 vccd1 vccd1 _14590_/C sky130_fd_sc_hd__a21o_1
X_16327_ _16327_/CLK _16327_/D vssd1 vssd1 vccd1 vccd1 _16327_/Q sky130_fd_sc_hd__dfxtp_2
X_13539_ _13539_/A vssd1 vssd1 vccd1 vccd1 _16020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16258_ _16268_/CLK _16258_/D vssd1 vssd1 vccd1 vccd1 _16258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15209_ _16224_/CLK _15209_/D vssd1 vssd1 vccd1 vccd1 _15209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16189_ _16189_/CLK _16189_/D vssd1 vssd1 vccd1 vccd1 _16189_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07962_ _07963_/A _07963_/B _07963_/C vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__a21oi_4
XFILLER_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09701_ _15412_/Q _09700_/C _09467_/X vssd1 vssd1 vccd1 vccd1 _09702_/B sky130_fd_sc_hd__a21oi_1
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07893_ _07893_/A _07893_/B vssd1 vssd1 vccd1 vccd1 _08152_/B sky130_fd_sc_hd__xor2_4
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _15400_/Q _09862_/B _09638_/C vssd1 vssd1 vccd1 vccd1 _09632_/Y sky130_fd_sc_hd__nand3_1
XFILLER_83_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09563_ _15391_/Q _09733_/B _09565_/C vssd1 vssd1 vccd1 vccd1 _09563_/X sky130_fd_sc_hd__and3_1
XFILLER_55_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08514_ _15231_/Q _08522_/C _13847_/A vssd1 vssd1 vccd1 vccd1 _08514_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09494_ _09519_/A _09494_/B _09494_/C vssd1 vssd1 vccd1 vccd1 _09495_/A sky130_fd_sc_hd__and3_1
X_08445_ _08435_/Y _08437_/X _08444_/Y vssd1 vssd1 vccd1 vccd1 _08446_/B sky130_fd_sc_hd__o21a_1
XFILLER_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08376_ _14414_/A vssd1 vssd1 vccd1 vccd1 _14363_/A sky130_fd_sc_hd__buf_2
XFILLER_136_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12910_ _15914_/Q _13018_/B _12914_/C vssd1 vssd1 vccd1 vccd1 _12910_/Y sky130_fd_sc_hd__nand3_1
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13890_ _14261_/A vssd1 vssd1 vccd1 vccd1 _13950_/B sky130_fd_sc_hd__buf_2
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12841_ _12838_/X _12839_/Y _12840_/Y _12836_/C vssd1 vssd1 vccd1 vccd1 _12843_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15194_/Q _15560_/D vssd1 vssd1 vccd1 vccd1 _15560_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _15893_/Q _12778_/C _12654_/X vssd1 vssd1 vccd1 vccd1 _12774_/C sky130_fd_sc_hd__a21o_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14552_/A _14511_/B _14511_/C vssd1 vssd1 vccd1 vccd1 _14512_/A sky130_fd_sc_hd__and3_1
X_11723_ _11723_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11727_/C sky130_fd_sc_hd__nor2_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15224_/Q _15491_/D vssd1 vssd1 vccd1 vccd1 _15491_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14442_/A _14442_/B vssd1 vssd1 vccd1 vccd1 _14442_/Y sky130_fd_sc_hd__nor2_1
X_11654_ _11654_/A vssd1 vssd1 vccd1 vccd1 _15715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _10602_/X _10603_/Y _10604_/Y _10600_/C vssd1 vssd1 vccd1 vccd1 _10607_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14373_ _14328_/X _14372_/X _14366_/B _14240_/X vssd1 vssd1 vccd1 vccd1 _14374_/B
+ sky130_fd_sc_hd__a31o_1
X_11585_ _15705_/Q _11697_/B _11585_/C vssd1 vssd1 vccd1 vccd1 _11585_/Y sky130_fd_sc_hd__nand3_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16112_ _16114_/CLK _16112_/D vssd1 vssd1 vccd1 vccd1 _16112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13324_ _13324_/A _13324_/B _13324_/C vssd1 vssd1 vccd1 vccd1 _13325_/C sky130_fd_sc_hd__nand3_1
XFILLER_128_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10536_ _10537_/B _10537_/C _10537_/A vssd1 vssd1 vccd1 vccd1 _10538_/B sky130_fd_sc_hd__a21o_1
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16043_ _16052_/CLK _16043_/D vssd1 vssd1 vccd1 vccd1 _16043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13255_ _13408_/A _13255_/B _13255_/C vssd1 vssd1 vccd1 vccd1 _13257_/B sky130_fd_sc_hd__or3_1
X_10467_ _10467_/A vssd1 vssd1 vccd1 vccd1 _15529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ _12206_/A vssd1 vssd1 vccd1 vccd1 _15802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _13700_/A vssd1 vssd1 vccd1 vccd1 _13394_/B sky130_fd_sc_hd__clkbuf_2
X_10398_ _10398_/A _10398_/B vssd1 vssd1 vccd1 vccd1 _10401_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12137_ _12150_/C vssd1 vssd1 vccd1 vccd1 _12159_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12068_ _12068_/A _12072_/C vssd1 vssd1 vccd1 vccd1 _12068_/X sky130_fd_sc_hd__or2_1
XFILLER_37_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11019_ _11019_/A _11019_/B _11019_/C vssd1 vssd1 vccd1 vccd1 _11020_/A sky130_fd_sc_hd__and3_1
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15827_ _15845_/CLK _15827_/D vssd1 vssd1 vccd1 vccd1 _15827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15758_ _15794_/CLK _15758_/D vssd1 vssd1 vccd1 vccd1 _15758_/Q sky130_fd_sc_hd__dfxtp_1
X_14709_ _14709_/A _14709_/B _14709_/C vssd1 vssd1 vccd1 vccd1 _14710_/C sky130_fd_sc_hd__nand3_1
X_15689_ _15763_/CLK _15689_/D vssd1 vssd1 vccd1 vccd1 _15689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _08231_/A _08231_/B _08231_/C vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__a21oi_1
XFILLER_119_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08161_ _10700_/A _07939_/B _08160_/X vssd1 vssd1 vccd1 vccd1 _08171_/B sky130_fd_sc_hd__o21ai_4
XFILLER_118_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08092_ _15485_/Q vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__inv_2
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08994_ _15303_/Q _09165_/B _09001_/C vssd1 vssd1 vccd1 vccd1 _08994_/X sky130_fd_sc_hd__and3_1
XFILLER_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ _07945_/A spike_out[1] _08420_/C vssd1 vssd1 vccd1 vccd1 _07946_/C sky130_fd_sc_hd__nor3_1
XFILLER_29_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07876_ _16053_/Q vssd1 vssd1 vccd1 vccd1 _13777_/C sky130_fd_sc_hd__inv_2
XFILLER_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09615_ _15399_/Q _09784_/B _09615_/C vssd1 vssd1 vccd1 vccd1 _09615_/X sky130_fd_sc_hd__and3_1
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ _09577_/C vssd1 vssd1 vccd1 vccd1 _09585_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09477_ _09476_/B _09476_/C _09307_/X vssd1 vssd1 vccd1 vccd1 _09478_/C sky130_fd_sc_hd__o21ai_1
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08428_ _08436_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08428_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ _08359_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _08359_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11370_ _15671_/Q _11601_/B _11374_/C vssd1 vssd1 vccd1 vccd1 _11370_/Y sky130_fd_sc_hd__nand3_1
XFILLER_109_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _10317_/X _10319_/Y _10320_/Y _10315_/C vssd1 vssd1 vccd1 vccd1 _10323_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13040_ _13071_/C vssd1 vssd1 vccd1 vccd1 _13078_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10252_ _10252_/A vssd1 vssd1 vccd1 vccd1 _15497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10183_ _15487_/Q _10239_/B _10191_/C vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__and3_1
XFILLER_133_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14991_ _14984_/B _14985_/C hold33/A _14989_/Y vssd1 vssd1 vccd1 vccd1 _14997_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13942_ _13942_/A _13942_/B _13942_/C vssd1 vssd1 vccd1 vccd1 _13943_/C sky130_fd_sc_hd__nand3_1
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13873_ _14379_/A vssd1 vssd1 vccd1 vccd1 _14117_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15612_ _15194_/Q _15612_/D vssd1 vssd1 vccd1 vccd1 _15612_/Q sky130_fd_sc_hd__dfxtp_2
X_12824_ _15901_/Q _12879_/B _12832_/C vssd1 vssd1 vccd1 vccd1 _12829_/A sky130_fd_sc_hd__and3_1
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15543_ _15655_/CLK _15543_/D vssd1 vssd1 vccd1 vccd1 _15543_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12755_ _13029_/A vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11702_/X _11703_/Y _11705_/Y _11700_/C vssd1 vssd1 vccd1 vccd1 _11708_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _15484_/CLK _15474_/D vssd1 vssd1 vccd1 vccd1 _15474_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _15878_/Q _12744_/B _12690_/C vssd1 vssd1 vccd1 vccd1 _12686_/Y sky130_fd_sc_hd__nand3_1
X_14425_ _16192_/Q _14447_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14427_/B sky130_fd_sc_hd__a21oi_1
X_11637_ _11635_/X _11636_/Y _11631_/B _11632_/C vssd1 vssd1 vccd1 vccd1 _11639_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14356_ _14353_/B _14352_/Y _14353_/A vssd1 vssd1 vccd1 vccd1 _14356_/Y sky130_fd_sc_hd__o21bai_1
X_11568_ _11661_/A _11568_/B _11573_/A vssd1 vssd1 vccd1 vccd1 _15702_/D sky130_fd_sc_hd__nor3_1
X_13307_ _13339_/A _13307_/B _13307_/C vssd1 vssd1 vccd1 vccd1 _13308_/A sky130_fd_sc_hd__and3_1
X_10519_ _10693_/A vssd1 vssd1 vccd1 vccd1 _10559_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14287_ _14287_/A vssd1 vssd1 vccd1 vccd1 _14287_/X sky130_fd_sc_hd__buf_2
X_11499_ _11538_/A _11499_/B _11499_/C vssd1 vssd1 vccd1 vccd1 _11500_/A sky130_fd_sc_hd__and3_1
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _16052_/CLK _16026_/D vssd1 vssd1 vccd1 vccd1 _16026_/Q sky130_fd_sc_hd__dfxtp_1
X_13238_ _13238_/A vssd1 vssd1 vccd1 vccd1 _15967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13169_ _13169_/A _13169_/B _13169_/C vssd1 vssd1 vccd1 vccd1 _13170_/C sky130_fd_sc_hd__nand3_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07730_ _15972_/Q _08132_/B vssd1 vssd1 vccd1 vccd1 _07740_/A sky130_fd_sc_hd__xnor2_4
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07661_ _12668_/A vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__clkbuf_4
X_09400_ _09398_/Y _09394_/C _09396_/X _09397_/Y vssd1 vssd1 vccd1 vccd1 _09401_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ _09331_/A vssd1 vssd1 vccd1 vccd1 _15354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ _09353_/A _09262_/B _09266_/A vssd1 vssd1 vccd1 vccd1 _15343_/D sky130_fd_sc_hd__nor3_1
X_08213_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08217_/A sky130_fd_sc_hd__xnor2_2
X_09193_ _09193_/A vssd1 vssd1 vccd1 vccd1 _15332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08144_ _15440_/Q _08144_/B vssd1 vssd1 vccd1 vccd1 _08144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08075_ _08075_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08305_/B sky130_fd_sc_hd__xnor2_1
XFILLER_106_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_130_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08977_ _08999_/A _08977_/B _08977_/C vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__and3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__buf_2
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_07928_ _07928_/A _07928_/B vssd1 vssd1 vccd1 vccd1 _07929_/B sky130_fd_sc_hd__nand2_2
XFILLER_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07859_ _12193_/A _07859_/B vssd1 vssd1 vccd1 vccd1 _07860_/B sky130_fd_sc_hd__nand2_1
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10870_ _10890_/C vssd1 vssd1 vccd1 vccd1 _10904_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09529_ _15385_/Q _09528_/C _09467_/X vssd1 vssd1 vccd1 vccd1 _09530_/B sky130_fd_sc_hd__a21oi_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12540_ _15857_/Q _12653_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12543_/B sky130_fd_sc_hd__nand3_1
XFILLER_61_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12471_ _12583_/A _12471_/B _12471_/C vssd1 vssd1 vccd1 vccd1 _12474_/B sky130_fd_sc_hd__or3_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14210_ _16148_/Q _14216_/C _13982_/X vssd1 vssd1 vccd1 vccd1 _14212_/C sky130_fd_sc_hd__a21o_1
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11422_ _11422_/A vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__clkbuf_2
X_15190_ _13920_/A _15188_/A _08335_/X vssd1 vssd1 vccd1 vccd1 _15191_/B sky130_fd_sc_hd__o21ai_1
XFILLER_137_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14141_ _14136_/Y _14139_/X _14140_/Y vssd1 vssd1 vccd1 vccd1 _16130_/D sky130_fd_sc_hd__o21a_1
X_11353_ _15670_/Q _11525_/B _11355_/C vssd1 vssd1 vccd1 vccd1 _11353_/X sky130_fd_sc_hd__and3_1
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _15507_/Q _10363_/B _10304_/C vssd1 vssd1 vccd1 vccd1 _10304_/X sky130_fd_sc_hd__and3_1
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ _14098_/A _14072_/B _14077_/A vssd1 vssd1 vccd1 vccd1 _16117_/D sky130_fd_sc_hd__nor3_1
X_11284_ _15659_/Q _11289_/C _11222_/X vssd1 vssd1 vccd1 vccd1 _11286_/C sky130_fd_sc_hd__a21o_1
XFILLER_106_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13023_ _15934_/Q _13022_/C _10970_/C vssd1 vssd1 vccd1 vccd1 _13024_/B sky130_fd_sc_hd__a21oi_1
X_10235_ _10247_/C vssd1 vssd1 vccd1 vccd1 _10256_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10166_ _10166_/A _10166_/B vssd1 vssd1 vccd1 vccd1 _10171_/C sky130_fd_sc_hd__nor2_1
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10097_ _10097_/A _10097_/B _10097_/C vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__and3_1
X_14974_ _16305_/Q vssd1 vssd1 vccd1 vccd1 _14981_/C sky130_fd_sc_hd__inv_2
XFILLER_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _14325_/A vssd1 vssd1 vccd1 vccd1 _13925_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13856_ _13856_/A _13856_/B vssd1 vssd1 vccd1 vccd1 _13857_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12807_ _12813_/B _12807_/B vssd1 vssd1 vccd1 vccd1 _12809_/A sky130_fd_sc_hd__or2_1
X_13787_ _13785_/X _13786_/Y _13782_/B _13783_/C vssd1 vssd1 vccd1 vccd1 _13789_/B
+ sky130_fd_sc_hd__o211ai_1
X_10999_ _15615_/Q _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__and3_1
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15526_ _15655_/CLK _15526_/D vssd1 vssd1 vccd1 vccd1 _15526_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12735_/X _12736_/Y _12737_/Y _12732_/C vssd1 vssd1 vccd1 vccd1 _12740_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15457_ _15484_/CLK _15457_/D vssd1 vssd1 vccd1 vccd1 _15457_/Q sky130_fd_sc_hd__dfxtp_1
X_12669_ _15877_/Q _12670_/C _12668_/X vssd1 vssd1 vccd1 vccd1 _12669_/Y sky130_fd_sc_hd__a21oi_1
X_14408_ _14408_/A vssd1 vssd1 vccd1 vccd1 _14408_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15388_ _15484_/CLK _15388_/D vssd1 vssd1 vccd1 vccd1 _15388_/Q sky130_fd_sc_hd__dfxtp_1
X_14339_ _16175_/Q _14468_/B _14345_/C vssd1 vssd1 vccd1 vccd1 _14342_/B sky130_fd_sc_hd__nand3_1
XFILLER_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08900_ _08900_/A vssd1 vssd1 vccd1 vccd1 _15287_/D sky130_fd_sc_hd__clkbuf_1
X_16009_ _16011_/CLK _16009_/D vssd1 vssd1 vccd1 vccd1 _16009_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09880_ _09878_/A _09878_/B _09879_/X vssd1 vssd1 vccd1 vccd1 _15438_/D sky130_fd_sc_hd__a21oi_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _15278_/Q _09067_/B _08831_/C vssd1 vssd1 vccd1 vccd1 _08839_/B sky130_fd_sc_hd__and3_1
XFILLER_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _15266_/Q _08996_/B _08769_/C vssd1 vssd1 vccd1 vccd1 _08762_/Y sky130_fd_sc_hd__nand3_1
XFILLER_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07713_ _07710_/X _07703_/A _15175_/A vssd1 vssd1 vccd1 vccd1 _07713_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08693_ _15257_/Q _08694_/C _08634_/X vssd1 vssd1 vccd1 vccd1 _08693_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07644_ _14300_/A vssd1 vssd1 vccd1 vccd1 _14634_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09314_ _09334_/C vssd1 vssd1 vccd1 vccd1 _09348_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09245_ _09245_/A _09245_/B vssd1 vssd1 vccd1 vccd1 _09247_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09176_ _09183_/A _09174_/Y _09175_/Y _09171_/C vssd1 vssd1 vccd1 vccd1 _09178_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ _08127_/A vssd1 vssd1 vccd1 vccd1 _15165_/C sky130_fd_sc_hd__buf_2
XFILLER_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08058_ _08058_/A vssd1 vssd1 vccd1 vccd1 _08062_/A sky130_fd_sc_hd__inv_2
XFILLER_134_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10020_ _10035_/A _10020_/B _10020_/C vssd1 vssd1 vccd1 vccd1 _10021_/A sky130_fd_sc_hd__and3_1
XFILLER_102_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11971_ _12084_/A _11971_/B _11975_/A vssd1 vssd1 vccd1 vccd1 _15765_/D sky130_fd_sc_hd__nor3_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13710_ _13716_/B _13710_/B vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__or2_1
X_10922_ _10960_/A _10922_/B _10922_/C vssd1 vssd1 vccd1 vccd1 _10923_/A sky130_fd_sc_hd__and3_1
XFILLER_44_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14690_ _07688_/X _14693_/C _07690_/X vssd1 vssd1 vccd1 vccd1 _14691_/B sky130_fd_sc_hd__o21ai_1
XFILLER_112_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _16041_/Q _13838_/B _13648_/C vssd1 vssd1 vccd1 vccd1 _13641_/X sky130_fd_sc_hd__and3_1
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10853_ _10931_/A _10853_/B _10858_/B vssd1 vssd1 vccd1 vccd1 _15590_/D sky130_fd_sc_hd__nor3_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16364_/CLK _16360_/D vssd1 vssd1 vccd1 vccd1 _16360_/Q sky130_fd_sc_hd__dfxtp_2
X_13572_ _13597_/C vssd1 vssd1 vccd1 vccd1 _13605_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10784_ _15581_/Q _10792_/C _10610_/X vssd1 vssd1 vccd1 vccd1 _10784_/Y sky130_fd_sc_hd__a21oi_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15311_ _15312_/CLK _15311_/D vssd1 vssd1 vccd1 vccd1 _15311_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12523_/A _12523_/B vssd1 vssd1 vccd1 vccd1 _12527_/C sky130_fd_sc_hd__nor2_1
X_16291_ _16304_/CLK _16291_/D vssd1 vssd1 vccd1 vccd1 _16291_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _15259_/CLK _15242_/D vssd1 vssd1 vccd1 vccd1 _15242_/Q sky130_fd_sc_hd__dfxtp_1
X_12454_ _12454_/A _12454_/B _12454_/C vssd1 vssd1 vccd1 vccd1 _12455_/A sky130_fd_sc_hd__and3_1
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11405_ _11420_/A _11405_/B _11405_/C vssd1 vssd1 vccd1 vccd1 _11406_/A sky130_fd_sc_hd__and3_1
XFILLER_138_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15173_ _15179_/A _15172_/Y _15168_/B _15169_/C vssd1 vssd1 vccd1 vccd1 _15175_/B
+ sky130_fd_sc_hd__o211a_1
X_12385_ _15832_/Q _12386_/C _12384_/X vssd1 vssd1 vccd1 vccd1 _12385_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_125_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14124_ _14124_/A vssd1 vssd1 vccd1 vccd1 _16127_/D sky130_fd_sc_hd__clkbuf_1
X_11336_ _11624_/A vssd1 vssd1 vccd1 vccd1 _11336_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_98_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14055_ _13912_/X _14053_/B _14054_/Y vssd1 vssd1 vccd1 vccd1 _16113_/D sky130_fd_sc_hd__o21a_1
X_11267_ _11267_/A vssd1 vssd1 vccd1 vccd1 _11309_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13006_ _13004_/Y _13000_/C _13002_/X _13003_/Y vssd1 vssd1 vccd1 vccd1 _13007_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10218_ _10216_/Y _10210_/C _10223_/A _10215_/Y vssd1 vssd1 vccd1 vccd1 _10223_/B
+ sky130_fd_sc_hd__a211oi_1
X_11198_ _15646_/Q _11431_/B _11198_/C vssd1 vssd1 vccd1 vccd1 _11208_/B sky130_fd_sc_hd__and3_1
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10149_ _15482_/Q _10155_/C _10030_/X vssd1 vssd1 vccd1 vccd1 _10149_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14957_ _14957_/A _14957_/B vssd1 vssd1 vccd1 vccd1 _14958_/B sky130_fd_sc_hd__nor2_1
XFILLER_94_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _13901_/Y _13906_/X _13907_/Y vssd1 vssd1 vccd1 vccd1 _16085_/D sky130_fd_sc_hd__o21a_1
X_14888_ _14766_/X _14891_/C _14808_/X vssd1 vssd1 vccd1 vccd1 _14889_/B sky130_fd_sc_hd__o21ai_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13839_ _16077_/Q _13846_/C _13693_/X vssd1 vssd1 vccd1 vccd1 _13839_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15509_ _15224_/Q _15509_/D vssd1 vssd1 vccd1 vccd1 _15509_/Q sky130_fd_sc_hd__dfxtp_1
X_09030_ _15308_/Q _09067_/C _09029_/X vssd1 vssd1 vccd1 vccd1 _09032_/B sky130_fd_sc_hd__a21oi_1
XFILLER_144_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09932_ _15448_/Q _09931_/C _09755_/X vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__a21oi_1
XFILLER_104_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09863_ _09860_/X _09861_/Y _09862_/Y _09858_/C vssd1 vssd1 vccd1 vccd1 _09865_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _08821_/A _08814_/B _08814_/C vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__and3_1
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _10663_/A vssd1 vssd1 vccd1 vccd1 _09794_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08745_ _15265_/Q _08919_/B _08745_/C vssd1 vssd1 vccd1 vccd1 _08745_/X sky130_fd_sc_hd__and3_1
XFILLER_66_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _15254_/Q _08715_/C _07623_/X vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__a21oi_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _08722_/A vssd1 vssd1 vccd1 vccd1 _15017_/A sky130_fd_sc_hd__buf_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ _15339_/Q _09451_/B _09236_/C vssd1 vssd1 vccd1 vccd1 _09228_/X sky130_fd_sc_hd__and3_1
XFILLER_127_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09159_ _15329_/Q _09160_/C _08929_/X vssd1 vssd1 vccd1 vccd1 _09159_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ _12170_/A _12170_/B _12170_/C vssd1 vssd1 vccd1 vccd1 _12171_/A sky130_fd_sc_hd__and3_1
XFILLER_135_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11121_ _15633_/Q _11121_/B _11121_/C vssd1 vssd1 vccd1 vccd1 _11121_/Y sky130_fd_sc_hd__nand3_1
XFILLER_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11052_ _15623_/Q _11058_/C _10933_/X vssd1 vssd1 vccd1 vccd1 _11054_/C sky130_fd_sc_hd__a21o_1
XFILLER_67_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10003_ _10016_/C vssd1 vssd1 vccd1 vccd1 _10024_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15860_ _15907_/CLK _15860_/D vssd1 vssd1 vccd1 vccd1 _15860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14811_ _14853_/A _14811_/B _14811_/C vssd1 vssd1 vccd1 vccd1 _14813_/A sky130_fd_sc_hd__and3_1
XFILLER_92_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15791_ _15809_/CLK _15791_/D vssd1 vssd1 vccd1 vccd1 _15791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11954_ _11954_/A _11954_/B vssd1 vssd1 vccd1 vccd1 _11958_/C sky130_fd_sc_hd__nor2_1
X_14742_ _14825_/A _14742_/B _14747_/A vssd1 vssd1 vccd1 vccd1 _16261_/D sky130_fd_sc_hd__nor3_1
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10905_ _15600_/Q _10910_/C _10848_/X vssd1 vssd1 vccd1 vccd1 _10905_/Y sky130_fd_sc_hd__a21oi_1
X_14673_ _16249_/Q _14677_/C _07649_/X vssd1 vssd1 vccd1 vccd1 _14673_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ _15753_/Q _11943_/B _11885_/C vssd1 vssd1 vccd1 vccd1 _11894_/A sky130_fd_sc_hd__and3_1
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13624_ _13648_/C vssd1 vssd1 vccd1 vccd1 _13655_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10836_ _10831_/X _10832_/Y _10835_/Y _10829_/C vssd1 vssd1 vccd1 vccd1 _10838_/B
+ sky130_fd_sc_hd__o211ai_1
Xrepeater11 _15196_/Q vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__buf_12
XFILLER_32_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16343_ _16344_/CLK _16343_/D vssd1 vssd1 vccd1 vccd1 _16343_/Q sky130_fd_sc_hd__dfxtp_2
X_13555_ _16025_/Q _13554_/C _13452_/X vssd1 vssd1 vccd1 vccd1 _13556_/B sky130_fd_sc_hd__a21oi_1
X_10767_ _10767_/A _10767_/B _10767_/C vssd1 vssd1 vccd1 vccd1 _10768_/C sky130_fd_sc_hd__nand3_1
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _15851_/Q _12512_/C _12332_/X vssd1 vssd1 vccd1 vccd1 _12506_/Y sky130_fd_sc_hd__a21oi_1
X_16274_ _16283_/CLK _16274_/D vssd1 vssd1 vccd1 vccd1 _16274_/Q sky130_fd_sc_hd__dfxtp_1
X_13486_ _13484_/X _13485_/Y _13480_/B _13481_/C vssd1 vssd1 vccd1 vccd1 _13488_/B
+ sky130_fd_sc_hd__o211ai_1
X_10698_ _10983_/A vssd1 vssd1 vccd1 vccd1 _10698_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15225_ _15259_/CLK _15225_/D vssd1 vssd1 vccd1 vccd1 _15225_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12437_ _12431_/B _12432_/C _12434_/X _12435_/Y vssd1 vssd1 vccd1 vccd1 _12438_/C
+ sky130_fd_sc_hd__a211o_1
X_15156_ _13920_/A _15154_/A _15086_/X vssd1 vssd1 vccd1 vccd1 _15157_/B sky130_fd_sc_hd__o21ai_1
X_12368_ _12368_/A _12368_/B _12373_/A vssd1 vssd1 vccd1 vccd1 _15828_/D sky130_fd_sc_hd__nor3_1
XFILLER_5_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _14106_/B _14106_/C _13919_/A vssd1 vssd1 vccd1 vccd1 _14108_/C sky130_fd_sc_hd__o21ai_1
X_11319_ _11326_/B _11319_/B vssd1 vssd1 vccd1 vccd1 _11321_/A sky130_fd_sc_hd__or2_1
XFILLER_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15087_ _13920_/A _15084_/A _15086_/X vssd1 vssd1 vccd1 vccd1 _15088_/B sky130_fd_sc_hd__o21ai_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12299_ _12299_/A _12299_/B _12299_/C vssd1 vssd1 vccd1 vccd1 _12301_/B sky130_fd_sc_hd__or3_1
X_14038_ _16114_/Q _14221_/B _14046_/C vssd1 vssd1 vccd1 vccd1 _14041_/A sky130_fd_sc_hd__and3_1
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15989_ _16052_/CLK _15989_/D vssd1 vssd1 vccd1 vccd1 _15989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08530_ input7/X vssd1 vssd1 vccd1 vccd1 _09699_/A sky130_fd_sc_hd__buf_2
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08461_ _08446_/A _08446_/B _08453_/B _08453_/A _08443_/A vssd1 vssd1 vccd1 vccd1
+ _08465_/C sky130_fd_sc_hd__o221a_1
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08392_ _08368_/A _08368_/B _08391_/X vssd1 vssd1 vccd1 vccd1 _08393_/B sky130_fd_sc_hd__a21o_2
XFILLER_149_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ _09185_/A _09018_/C vssd1 vssd1 vccd1 vccd1 _09013_/X sky130_fd_sc_hd__or2_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09915_ _09915_/A vssd1 vssd1 vccd1 vccd1 _15444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09846_ _10134_/A vssd1 vssd1 vccd1 vccd1 _10074_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09777_ _15425_/Q _10010_/B _09784_/C vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__nand3_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08728_ _08765_/A _08728_/B _08728_/C vssd1 vssd1 vccd1 vccd1 _08729_/A sky130_fd_sc_hd__and3_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08667_/B _08659_/B vssd1 vssd1 vccd1 vccd1 _08663_/A sky130_fd_sc_hd__or2_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11727_/A _11670_/B _11670_/C vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__or3_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10621_ _10619_/Y _10615_/C _10627_/A _10618_/Y vssd1 vssd1 vccd1 vccd1 _10627_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13340_ _13340_/A vssd1 vssd1 vccd1 vccd1 _15985_/D sky130_fd_sc_hd__clkbuf_1
X_10552_ _10559_/A _10552_/B _10552_/C vssd1 vssd1 vccd1 vccd1 _10553_/A sky130_fd_sc_hd__and3_1
XFILLER_139_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13271_ _13272_/B _13272_/C _13272_/A vssd1 vssd1 vccd1 vccd1 _13273_/B sky130_fd_sc_hd__a21o_1
XFILLER_139_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10483_ _10483_/A vssd1 vssd1 vccd1 vccd1 _15532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15010_ _15051_/A _15010_/B _15010_/C vssd1 vssd1 vccd1 vccd1 _15012_/A sky130_fd_sc_hd__and3_1
X_12222_ _15806_/Q _12228_/C _12048_/X vssd1 vssd1 vccd1 vccd1 _12222_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12153_ _12147_/B _12148_/C _12150_/X _12151_/Y vssd1 vssd1 vccd1 vccd1 _12154_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _15631_/Q _11143_/C _11047_/X vssd1 vssd1 vccd1 vccd1 _11106_/B sky130_fd_sc_hd__a21oi_1
X_12084_ _12084_/A _12084_/B _12089_/A vssd1 vssd1 vccd1 vccd1 _15783_/D sky130_fd_sc_hd__nor3_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11035_ _11267_/A vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15912_ _07603_/A _15912_/D vssd1 vssd1 vccd1 vccd1 _15912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15843_ _15907_/CLK _15843_/D vssd1 vssd1 vccd1 vccd1 _15843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15774_ _15794_/CLK _15774_/D vssd1 vssd1 vccd1 vccd1 _15774_/Q sky130_fd_sc_hd__dfxtp_2
X_12986_ _13016_/C vssd1 vssd1 vccd1 vccd1 _13022_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14725_ _14720_/A _14723_/B _14646_/X vssd1 vssd1 vccd1 vccd1 _14731_/C sky130_fd_sc_hd__o21a_1
X_11937_ _15761_/Q _11943_/C _11760_/X vssd1 vssd1 vccd1 vccd1 _11937_/Y sky130_fd_sc_hd__a21oi_1
X_11868_ _11868_/A vssd1 vssd1 vccd1 vccd1 _15749_/D sky130_fd_sc_hd__clkbuf_1
X_14656_ _14656_/A _14656_/B vssd1 vssd1 vccd1 vccd1 _16240_/D sky130_fd_sc_hd__nor2_1
XFILLER_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10819_ _15587_/Q _10876_/B _10825_/C vssd1 vssd1 vccd1 vccd1 _10822_/B sky130_fd_sc_hd__nand3_1
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13607_ _13613_/B _13607_/B vssd1 vssd1 vccd1 vccd1 _13609_/A sky130_fd_sc_hd__or2_1
X_11799_ _15740_/Q _11804_/C _11798_/X vssd1 vssd1 vccd1 vccd1 _11801_/C sky130_fd_sc_hd__a21o_1
X_14587_ _16229_/Q _14587_/B _14593_/C vssd1 vssd1 vccd1 vccd1 _14590_/B sky130_fd_sc_hd__nand3_1
X_16326_ _16344_/CLK _16326_/D vssd1 vssd1 vccd1 vccd1 _16326_/Q sky130_fd_sc_hd__dfxtp_2
X_13538_ _13538_/A _13538_/B _13538_/C vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__and3_1
X_16257_ _16268_/CLK _16257_/D vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
X_13469_ _15999_/Q vssd1 vssd1 vccd1 vccd1 _13475_/C sky130_fd_sc_hd__inv_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15208_ _16353_/CLK _15208_/D vssd1 vssd1 vccd1 vccd1 _15208_/Q sky130_fd_sc_hd__dfxtp_1
X_16188_ _16204_/CLK _16188_/D vssd1 vssd1 vccd1 vccd1 _16188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15139_ _15145_/A _15138_/Y _15134_/B _15135_/C vssd1 vssd1 vccd1 vccd1 _15141_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07961_ _15061_/C _07917_/B _07916_/A vssd1 vssd1 vccd1 vccd1 _07963_/C sky130_fd_sc_hd__o21a_1
XFILLER_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _15412_/Q _09931_/B _09700_/C vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__and3_1
X_07892_ _09658_/A _07892_/B vssd1 vssd1 vccd1 vccd1 _07893_/B sky130_fd_sc_hd__xnor2_2
XFILLER_68_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09631_ _10785_/A vssd1 vssd1 vccd1 vccd1 _09862_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09562_ _09562_/A vssd1 vssd1 vccd1 vccd1 _15389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08513_ _12616_/A vssd1 vssd1 vccd1 vccd1 _13847_/A sky130_fd_sc_hd__buf_4
XFILLER_82_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09493_ _09493_/A _09493_/B _09493_/C vssd1 vssd1 vccd1 vccd1 _09494_/C sky130_fd_sc_hd__nand3_1
XFILLER_36_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08444_ _08444_/A _08444_/B vssd1 vssd1 vccd1 vccd1 _08444_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08375_ _08375_/A _08375_/B vssd1 vssd1 vccd1 vccd1 _08378_/A sky130_fd_sc_hd__or2_1
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09829_ _09829_/A vssd1 vssd1 vccd1 vccd1 _15430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12840_ _15903_/Q _12840_/B _12840_/C vssd1 vssd1 vccd1 vccd1 _12840_/Y sky130_fd_sc_hd__nand3_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12771_ _15893_/Q _12935_/B _12778_/C vssd1 vssd1 vccd1 vccd1 _12774_/B sky130_fd_sc_hd__nand3_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11722_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__nor2_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _14510_/A _14510_/B _14510_/C vssd1 vssd1 vccd1 vccd1 _14511_/C sky130_fd_sc_hd__nand3_1
X_15490_ _15224_/Q _15490_/D vssd1 vssd1 vccd1 vccd1 _15490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11653_ _11653_/A _11653_/B _11653_/C vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__and3_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _16195_/Q _14447_/C _14395_/X vssd1 vssd1 vccd1 vccd1 _14443_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10604_ _15552_/Q _10778_/B _10604_/C vssd1 vssd1 vccd1 vccd1 _10604_/Y sky130_fd_sc_hd__nand3_1
X_14372_ _14372_/A vssd1 vssd1 vccd1 vccd1 _14372_/X sky130_fd_sc_hd__clkbuf_2
X_11584_ _15706_/Q _11585_/C _11526_/X vssd1 vssd1 vccd1 vccd1 _11584_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ _13324_/B _13324_/C _13324_/A vssd1 vssd1 vccd1 vccd1 _13325_/B sky130_fd_sc_hd__a21o_1
X_16111_ _16114_/CLK _16111_/D vssd1 vssd1 vccd1 vccd1 _16111_/Q sky130_fd_sc_hd__dfxtp_1
X_10535_ _15542_/Q _10540_/C _10357_/X vssd1 vssd1 vccd1 vccd1 _10537_/C sky130_fd_sc_hd__a21o_1
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13254_ _13252_/A _13252_/B _13253_/X vssd1 vssd1 vccd1 vccd1 _15969_/D sky130_fd_sc_hd__a21oi_1
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16042_ _16052_/CLK _16042_/D vssd1 vssd1 vccd1 vccd1 _16042_/Q sky130_fd_sc_hd__dfxtp_1
X_10466_ _10503_/A _10466_/B _10466_/C vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__and3_1
X_12205_ _12226_/A _12205_/B _12205_/C vssd1 vssd1 vccd1 vccd1 _12206_/A sky130_fd_sc_hd__and3_1
XFILLER_136_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _13185_/A vssd1 vssd1 vccd1 vccd1 _15958_/D sky130_fd_sc_hd__clkbuf_1
X_10397_ _10405_/B _10397_/B vssd1 vssd1 vccd1 vccd1 _10401_/A sky130_fd_sc_hd__or2_1
XFILLER_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12136_ _15791_/Q vssd1 vssd1 vccd1 vccd1 _12150_/C sky130_fd_sc_hd__inv_2
XFILLER_145_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12067_ _12067_/A _12067_/B vssd1 vssd1 vccd1 vccd1 _12072_/C sky130_fd_sc_hd__nor2_1
X_11018_ _11016_/Y _11011_/C _11014_/X _11015_/Y vssd1 vssd1 vccd1 vccd1 _11019_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15826_ _15907_/CLK _15826_/D vssd1 vssd1 vccd1 vccd1 _15826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15757_ _15794_/CLK _15757_/D vssd1 vssd1 vccd1 vccd1 _15757_/Q sky130_fd_sc_hd__dfxtp_1
X_12969_ _15925_/Q _12968_/C _10970_/C vssd1 vssd1 vccd1 vccd1 _12970_/B sky130_fd_sc_hd__a21oi_1
XFILLER_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14708_ _14709_/B _14709_/C _14709_/A vssd1 vssd1 vccd1 vccd1 _14710_/B sky130_fd_sc_hd__a21o_1
X_15688_ _15763_/CLK _15688_/D vssd1 vssd1 vccd1 vccd1 _15688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14639_ hold26/A _14755_/B _14639_/C vssd1 vssd1 vccd1 vccd1 _14641_/A sky130_fd_sc_hd__and3_1
XFILLER_14_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08160_ _08731_/A _08160_/B vssd1 vssd1 vccd1 vccd1 _08160_/X sky130_fd_sc_hd__or2_1
X_16309_ _16312_/CLK _16309_/D vssd1 vssd1 vccd1 vccd1 _16309_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ _15503_/Q vssd1 vssd1 vccd1 vccd1 _10289_/A sky130_fd_sc_hd__inv_2
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08993_ _08993_/A vssd1 vssd1 vccd1 vccd1 _15301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07944_ _07945_/A spike_out[1] _08420_/C vssd1 vssd1 vccd1 vccd1 _07946_/B sky130_fd_sc_hd__o21a_1
XFILLER_87_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07875_ _16080_/Q vssd1 vssd1 vccd1 vccd1 _13937_/C sky130_fd_sc_hd__clkinv_2
XFILLER_110_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09614_ _09614_/A vssd1 vssd1 vccd1 vccd1 _15397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _09565_/C vssd1 vssd1 vccd1 vccd1 _09577_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09476_ _09708_/A _09476_/B _09476_/C vssd1 vssd1 vccd1 vccd1 _09478_/B sky130_fd_sc_hd__or3_1
XFILLER_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08427_ state1[3] _08433_/A vssd1 vssd1 vccd1 vccd1 _08436_/B sky130_fd_sc_hd__and2_1
X_08358_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__xnor2_2
XFILLER_109_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08289_ _08289_/A _08221_/A vssd1 vssd1 vccd1 vccd1 _08289_/X sky130_fd_sc_hd__or2b_1
XFILLER_137_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ _15508_/Q _10441_/B _10325_/C vssd1 vssd1 vccd1 vccd1 _10320_/Y sky130_fd_sc_hd__nand3_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10251_ _10266_/A _10251_/B _10251_/C vssd1 vssd1 vccd1 vccd1 _10252_/A sky130_fd_sc_hd__and3_1
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10182_ _15487_/Q _10220_/C _10181_/X vssd1 vssd1 vccd1 vccd1 _10184_/B sky130_fd_sc_hd__a21oi_1
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14990_ hold33/A _14989_/Y _14984_/B _14985_/C vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__o211a_1
XFILLER_93_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13941_ _13942_/B _13942_/C _13942_/A vssd1 vssd1 vccd1 vccd1 _13943_/B sky130_fd_sc_hd__a21o_1
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13872_ _16084_/Q _13903_/C _13822_/X vssd1 vssd1 vccd1 vccd1 _13875_/B sky130_fd_sc_hd__a21oi_1
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15611_ _15620_/CLK _15611_/D vssd1 vssd1 vccd1 vccd1 _15611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12823_ _15901_/Q _12861_/C _12767_/X vssd1 vssd1 vccd1 vccd1 _12825_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15542_ _15655_/CLK _15542_/D vssd1 vssd1 vccd1 vccd1 _15542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12752_/A _12752_/B _12753_/X vssd1 vssd1 vccd1 vccd1 _15888_/D sky130_fd_sc_hd__a21oi_1
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _15724_/Q _11938_/B _11712_/C vssd1 vssd1 vccd1 vccd1 _11705_/Y sky130_fd_sc_hd__nand3_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15473_ _15483_/CLK _15473_/D vssd1 vssd1 vccd1 vccd1 _15473_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _15879_/Q _12690_/C _12569_/X vssd1 vssd1 vccd1 vccd1 _12685_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11636_ _15714_/Q _11643_/C _11519_/X vssd1 vssd1 vccd1 vccd1 _11636_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14424_ _14435_/C vssd1 vssd1 vccd1 vccd1 _14447_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14355_ _14353_/A _14353_/B _14352_/Y _14354_/Y vssd1 vssd1 vccd1 vccd1 _16174_/D
+ sky130_fd_sc_hd__o31a_1
X_11567_ _15703_/Q _11737_/B _11576_/C vssd1 vssd1 vccd1 vccd1 _11573_/A sky130_fd_sc_hd__and3_1
XFILLER_143_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10518_ _10516_/A _10516_/B _10517_/X vssd1 vssd1 vccd1 vccd1 _15537_/D sky130_fd_sc_hd__a21oi_1
X_13306_ _13304_/B _13304_/C _13305_/X vssd1 vssd1 vccd1 vccd1 _13307_/C sky130_fd_sc_hd__o21ai_1
X_14286_ _14299_/C vssd1 vssd1 vccd1 vccd1 _14313_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11498_ _11497_/B _11497_/C _11327_/X vssd1 vssd1 vccd1 vccd1 _11499_/C sky130_fd_sc_hd__o21ai_1
XFILLER_6_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13237_ _13281_/A _13237_/B _13237_/C vssd1 vssd1 vccd1 vccd1 _13238_/A sky130_fd_sc_hd__and3_1
X_16025_ _16052_/CLK _16025_/D vssd1 vssd1 vccd1 vccd1 _16025_/Q sky130_fd_sc_hd__dfxtp_1
X_10449_ _15527_/Q _10681_/B _10453_/C vssd1 vssd1 vccd1 vccd1 _10449_/Y sky130_fd_sc_hd__nand3_1
XFILLER_108_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13168_ _13169_/B _13169_/C _13169_/A vssd1 vssd1 vccd1 vccd1 _13170_/B sky130_fd_sc_hd__a21o_1
XFILLER_124_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12119_ _12117_/Y _12112_/C _12124_/A _12116_/Y vssd1 vssd1 vccd1 vccd1 _12124_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_111_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13099_ _13099_/A vssd1 vssd1 vccd1 vccd1 _13679_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ _10947_/A vssd1 vssd1 vccd1 vccd1 _12668_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15809_ _15809_/CLK _15809_/D vssd1 vssd1 vccd1 vccd1 _15809_/Q sky130_fd_sc_hd__dfxtp_1
X_09330_ _09345_/A _09330_/B _09330_/C vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__and3_1
XFILLER_34_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09261_ _15344_/Q _09372_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09266_/A sky130_fd_sc_hd__and3_1
XFILLER_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08212_ _08064_/A _08064_/B _08211_/Y vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__a21oi_2
X_09192_ _09233_/A _09192_/B _09192_/C vssd1 vssd1 vccd1 vccd1 _09193_/A sky130_fd_sc_hd__and3_1
X_08143_ _08143_/A _08143_/B vssd1 vssd1 vccd1 vccd1 _08260_/A sky130_fd_sc_hd__xnor2_4
XFILLER_147_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08074_ _08226_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_08976_ _08976_/A _08976_/B _08976_/C vssd1 vssd1 vccd1 vccd1 _08977_/C sky130_fd_sc_hd__nand3_1
Xhold25 hold8/X vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07927_ _15746_/Q _16341_/Q vssd1 vssd1 vccd1 vccd1 _07928_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07858_ _12193_/A _07859_/B vssd1 vssd1 vccd1 vccd1 _07860_/A sky130_fd_sc_hd__or2_1
XFILLER_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07789_ _15674_/Q vssd1 vssd1 vccd1 vccd1 _11388_/A sky130_fd_sc_hd__clkinv_4
XFILLER_37_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _15385_/Q _09644_/B _09528_/C vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__and3_1
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ _09459_/A vssd1 vssd1 vccd1 vccd1 _15373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12470_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12510_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11421_ _11421_/A vssd1 vssd1 vccd1 vccd1 _15679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14140_ _14136_/Y _14139_/X _14049_/X vssd1 vssd1 vccd1 vccd1 _14140_/Y sky130_fd_sc_hd__a21oi_1
X_11352_ _11352_/A vssd1 vssd1 vccd1 vccd1 _15668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10303_ _10303_/A vssd1 vssd1 vccd1 vccd1 _15505_/D sky130_fd_sc_hd__clkbuf_1
X_14071_ _16119_/Q _14071_/B _14071_/C vssd1 vssd1 vccd1 vccd1 _14077_/A sky130_fd_sc_hd__and3_1
X_11283_ _15659_/Q _11510_/B _11289_/C vssd1 vssd1 vccd1 vccd1 _11286_/B sky130_fd_sc_hd__nand3_1
X_13022_ _15934_/Q _13078_/B _13022_/C vssd1 vssd1 vccd1 vccd1 _13031_/B sky130_fd_sc_hd__and3_1
X_10234_ _10234_/A vssd1 vssd1 vccd1 vccd1 _10247_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10165_ _10165_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10166_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10096_ _10094_/Y _10088_/C _10092_/X _10093_/Y vssd1 vssd1 vccd1 vccd1 _10097_/C
+ sky130_fd_sc_hd__a211o_1
X_14973_ _16331_/Q _16330_/Q _16329_/Q _14818_/X vssd1 vssd1 vccd1 vccd1 _16314_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13924_ _13920_/X _13917_/B _13923_/Y vssd1 vssd1 vccd1 vccd1 _16087_/D sky130_fd_sc_hd__o21a_1
XFILLER_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13855_ _13861_/B _13855_/B vssd1 vssd1 vccd1 vccd1 _13857_/A sky130_fd_sc_hd__or2_1
X_12806_ _15898_/Q _12805_/C _12631_/X vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13786_ _16067_/Q _13785_/C _10950_/C vssd1 vssd1 vccd1 vccd1 _13786_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10998_ _10998_/A vssd1 vssd1 vccd1 vccd1 _15613_/D sky130_fd_sc_hd__clkbuf_1
X_15525_ _15655_/CLK _15525_/D vssd1 vssd1 vccd1 vccd1 _15525_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _15886_/Q _12793_/B _12742_/C vssd1 vssd1 vccd1 vccd1 _12737_/Y sky130_fd_sc_hd__nand3_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15456_ _15484_/CLK _15456_/D vssd1 vssd1 vccd1 vccd1 _15456_/Q sky130_fd_sc_hd__dfxtp_1
X_12668_ _12668_/A vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__buf_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14407_ _14401_/Y _14405_/X _14406_/Y vssd1 vssd1 vccd1 vccd1 _16184_/D sky130_fd_sc_hd__o21a_1
XFILLER_129_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ _15718_/Q _15717_/Q _15716_/Q _11560_/X vssd1 vssd1 vccd1 vccd1 _15710_/D
+ sky130_fd_sc_hd__o31a_1
X_15387_ _15484_/CLK _15387_/D vssd1 vssd1 vccd1 vccd1 _15387_/Q sky130_fd_sc_hd__dfxtp_2
X_12599_ _12621_/A _12599_/B _12599_/C vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__and3_1
XFILLER_128_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14338_ _14427_/A _14338_/B _14342_/A vssd1 vssd1 vccd1 vccd1 _16171_/D sky130_fd_sc_hd__nor3_1
XFILLER_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14269_ _16160_/Q _14357_/B _14269_/C vssd1 vssd1 vccd1 vccd1 _14269_/X sky130_fd_sc_hd__and3_1
X_16008_ _16031_/CLK _16008_/D vssd1 vssd1 vccd1 vccd1 _16008_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _09699_/A vssd1 vssd1 vccd1 vccd1 _09067_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _13693_/A vssd1 vssd1 vccd1 vccd1 _08996_/B sky130_fd_sc_hd__clkbuf_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07712_ _15181_/A vssd1 vssd1 vccd1 vccd1 _15175_/A sky130_fd_sc_hd__buf_2
X_08692_ _15257_/Q _08865_/B _08694_/C vssd1 vssd1 vccd1 vccd1 _08692_/X sky130_fd_sc_hd__and3_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07643_ _12609_/A vssd1 vssd1 vccd1 vccd1 _14300_/A sky130_fd_sc_hd__buf_4
XFILLER_81_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09313_ _09326_/C vssd1 vssd1 vccd1 vccd1 _09334_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16359_/CLK sky130_fd_sc_hd__clkbuf_16
X_09244_ _09251_/B _09244_/B vssd1 vssd1 vccd1 vccd1 _09247_/A sky130_fd_sc_hd__or2_1
X_09175_ _15330_/Q _09238_/B _09179_/C vssd1 vssd1 vccd1 vccd1 _09175_/Y sky130_fd_sc_hd__nand3_1
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08126_ _08546_/A _09024_/A _08125_/Y vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__o21ai_2
XFILLER_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08057_ _11562_/A _11676_/A _08056_/Y vssd1 vssd1 vccd1 vccd1 _08058_/A sky130_fd_sc_hd__o21ai_2
XFILLER_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08959_ _08957_/A _08957_/B _08958_/X vssd1 vssd1 vccd1 vccd1 _15295_/D sky130_fd_sc_hd__a21oi_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11970_ _15766_/Q _12025_/B _11978_/C vssd1 vssd1 vccd1 vccd1 _11975_/A sky130_fd_sc_hd__and3_1
XFILLER_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10921_ _10920_/B _10920_/C _10751_/X vssd1 vssd1 vccd1 vccd1 _10922_/C sky130_fd_sc_hd__o21ai_1
XFILLER_17_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10852_ _10850_/Y _10845_/C _10858_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _10858_/B
+ sky130_fd_sc_hd__a211oi_1
X_13640_ _13640_/A vssd1 vssd1 vccd1 vccd1 _13838_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _13583_/C vssd1 vssd1 vccd1 vccd1 _13597_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10783_ _15581_/Q _10895_/B _10792_/C vssd1 vssd1 vccd1 vccd1 _10783_/X sky130_fd_sc_hd__and3_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16241_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15310_ _15312_/CLK _15310_/D vssd1 vssd1 vccd1 vccd1 _15310_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12522_/A _12522_/B vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16304_/CLK _16290_/D vssd1 vssd1 vccd1 vccd1 _16290_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _15351_/CLK _15241_/D vssd1 vssd1 vccd1 vccd1 _15241_/Q sky130_fd_sc_hd__dfxtp_1
X_12453_ _12451_/Y _12446_/C _12449_/X _12450_/Y vssd1 vssd1 vccd1 vccd1 _12454_/C
+ sky130_fd_sc_hd__a211o_1
X_11404_ _11398_/B _11399_/C _11401_/X _11402_/Y vssd1 vssd1 vccd1 vccd1 _11405_/C
+ sky130_fd_sc_hd__a211o_1
X_12384_ _12668_/A vssd1 vssd1 vccd1 vccd1 _12384_/X sky130_fd_sc_hd__clkbuf_4
X_15172_ _16366_/Q _15176_/C _13286_/B vssd1 vssd1 vccd1 vccd1 _15172_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11335_ _11367_/C vssd1 vssd1 vccd1 vccd1 _11374_/C sky130_fd_sc_hd__clkbuf_2
X_14123_ _14123_/A _14123_/B _14123_/C vssd1 vssd1 vccd1 vccd1 _14124_/A sky130_fd_sc_hd__and3_1
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11266_ _11264_/A _11264_/B _11265_/X vssd1 vssd1 vccd1 vccd1 _15654_/D sky130_fd_sc_hd__a21oi_1
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14054_ _14054_/A _14054_/B vssd1 vssd1 vccd1 vccd1 _14054_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10217_ _10223_/A _10215_/Y _10216_/Y _10210_/C vssd1 vssd1 vccd1 vccd1 _10219_/B
+ sky130_fd_sc_hd__o211a_1
X_13005_ _13002_/X _13003_/Y _13004_/Y _13000_/C vssd1 vssd1 vccd1 vccd1 _13007_/B
+ sky130_fd_sc_hd__o211ai_1
X_11197_ _11197_/A vssd1 vssd1 vccd1 vccd1 _11431_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _15482_/Q _10317_/B _10155_/C vssd1 vssd1 vccd1 vccd1 _10148_/X sky130_fd_sc_hd__and3_1
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10079_ _10097_/A _10079_/B _10079_/C vssd1 vssd1 vccd1 vccd1 _10080_/A sky130_fd_sc_hd__and3_1
X_14956_ _14956_/A _14956_/B vssd1 vssd1 vccd1 vccd1 _14957_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13907_ _13901_/Y _13906_/X _08168_/X vssd1 vssd1 vccd1 vccd1 _13907_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14887_ _14963_/A _14891_/C vssd1 vssd1 vccd1 vccd1 _14889_/A sky130_fd_sc_hd__and2_1
X_13838_ _16077_/Q _13838_/B _13846_/C vssd1 vssd1 vccd1 vccd1 _13838_/X sky130_fd_sc_hd__and3_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13769_ _13769_/A vssd1 vssd1 vccd1 vccd1 _16060_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_42_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16187_/CLK sky130_fd_sc_hd__clkbuf_16
X_15508_ _15224_/Q _15508_/D vssd1 vssd1 vccd1 vccd1 _15508_/Q sky130_fd_sc_hd__dfxtp_1
X_15439_ _15484_/CLK _15439_/D vssd1 vssd1 vccd1 vccd1 _15439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _15448_/Q _09931_/B _09931_/C vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__and3_1
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09862_ _15436_/Q _09862_/B _09867_/C vssd1 vssd1 vccd1 vccd1 _09862_/Y sky130_fd_sc_hd__nand3_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08813_ _08811_/Y _08806_/C _08808_/X _08809_/Y vssd1 vssd1 vccd1 vccd1 _08814_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _15427_/Q _10022_/B _09796_/C vssd1 vssd1 vccd1 vccd1 _09793_/X sky130_fd_sc_hd__and3_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08744_ _08744_/A vssd1 vssd1 vccd1 vccd1 _15263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _08706_/C vssd1 vssd1 vccd1 vccd1 _08715_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_26_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _08421_/A _07626_/B _07638_/A vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__nor3_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16224_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09227_ _09801_/A vssd1 vssd1 vccd1 vccd1 _09451_/B sky130_fd_sc_hd__buf_2
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09158_ _15329_/Q _09158_/B _09160_/C vssd1 vssd1 vccd1 vccd1 _09158_/X sky130_fd_sc_hd__and3_1
XFILLER_135_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08109_ _08109_/A vssd1 vssd1 vccd1 vccd1 _15096_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09089_ _09202_/A _09089_/B _09093_/A vssd1 vssd1 vccd1 vccd1 _15316_/D sky130_fd_sc_hd__nor3_1
XFILLER_108_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11120_ _15634_/Q _11121_/C _10948_/X vssd1 vssd1 vccd1 vccd1 _11120_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _15623_/Q _11221_/B _11058_/C vssd1 vssd1 vccd1 vccd1 _11054_/B sky130_fd_sc_hd__nand3_1
XFILLER_107_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10002_ _10002_/A vssd1 vssd1 vccd1 vccd1 _10016_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14810_ _14810_/A _14810_/B vssd1 vssd1 vccd1 vccd1 _16275_/D sky130_fd_sc_hd__nor2_1
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15790_ _15195_/Q _15790_/D vssd1 vssd1 vccd1 vccd1 _15790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14741_ _16265_/Q _14778_/B _14743_/C vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__and3_1
X_11953_ _11953_/A _11953_/B vssd1 vssd1 vccd1 vccd1 _11954_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10904_ _15600_/Q _11078_/B _10904_/C vssd1 vssd1 vccd1 vccd1 _10914_/A sky130_fd_sc_hd__and3_1
XFILLER_72_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14672_ _16249_/Q _14833_/B _14677_/C vssd1 vssd1 vccd1 vccd1 _14680_/A sky130_fd_sc_hd__and3_1
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11884_ _11884_/A vssd1 vssd1 vccd1 vccd1 _15751_/D sky130_fd_sc_hd__clkbuf_1
X_13623_ _13634_/C vssd1 vssd1 vccd1 vccd1 _13648_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_10835_ _15588_/Q _11121_/B _10835_/C vssd1 vssd1 vccd1 vccd1 _10835_/Y sky130_fd_sc_hd__nand3_1
Xrepeater12 _15794_/CLK vssd1 vssd1 vccd1 vccd1 _15763_/CLK sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_24_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _16143_/CLK sky130_fd_sc_hd__clkbuf_16
X_16342_ _16352_/CLK _16342_/D vssd1 vssd1 vccd1 vccd1 _16342_/Q sky130_fd_sc_hd__dfxtp_2
X_13554_ _16025_/Q _13605_/B _13554_/C vssd1 vssd1 vccd1 vccd1 _13561_/B sky130_fd_sc_hd__and3_1
XFILLER_9_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10766_ _10767_/B _10767_/C _10767_/A vssd1 vssd1 vccd1 vccd1 _10768_/B sky130_fd_sc_hd__a21o_1
XFILLER_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12505_ _15851_/Q _12675_/B _12512_/C vssd1 vssd1 vccd1 vccd1 _12505_/X sky130_fd_sc_hd__and3_1
X_16273_ _16273_/CLK _16273_/D vssd1 vssd1 vccd1 vccd1 _16273_/Q sky130_fd_sc_hd__dfxtp_2
X_10697_ _10697_/A vssd1 vssd1 vccd1 vccd1 _15565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13485_ _16013_/Q _13484_/C _13277_/X vssd1 vssd1 vccd1 vccd1 _13485_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_145_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ _15485_/CLK _15224_/D vssd1 vssd1 vccd1 vccd1 _15224_/Q sky130_fd_sc_hd__dfxtp_4
X_12436_ _12434_/X _12435_/Y _12431_/B _12432_/C vssd1 vssd1 vccd1 vccd1 _12438_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_126_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15155_ _15189_/A _15189_/B _15155_/C vssd1 vssd1 vccd1 vccd1 _15157_/A sky130_fd_sc_hd__and3_1
X_12367_ _15829_/Q _12593_/B _12376_/C vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__and3_1
X_14106_ _14106_/A _14106_/B _14106_/C vssd1 vssd1 vccd1 vccd1 _14108_/B sky130_fd_sc_hd__or3_1
X_11318_ _15664_/Q _11317_/C _11199_/X vssd1 vssd1 vccd1 vccd1 _11319_/B sky130_fd_sc_hd__a21oi_1
XFILLER_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12298_ _12413_/A vssd1 vssd1 vccd1 vccd1 _12337_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15086_ _15086_/A vssd1 vssd1 vccd1 vccd1 _15086_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11249_ _11249_/A _11249_/B _11249_/C vssd1 vssd1 vccd1 vccd1 _11250_/A sky130_fd_sc_hd__and3_1
X_14037_ _14098_/A _14037_/B _14040_/B vssd1 vssd1 vccd1 vccd1 _16110_/D sky130_fd_sc_hd__nor3_1
XFILLER_141_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15988_ _16052_/CLK _15988_/D vssd1 vssd1 vccd1 vccd1 _15988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14939_ _16310_/Q _14977_/B _14941_/C vssd1 vssd1 vccd1 vccd1 _14945_/A sky130_fd_sc_hd__and3_1
X_08460_ _13972_/A vssd1 vssd1 vccd1 vccd1 _08519_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08391_ _08391_/A _08391_/B vssd1 vssd1 vccd1 vccd1 _08391_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_15_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _16031_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09012_ _09012_/A _09012_/B vssd1 vssd1 vccd1 vccd1 _09018_/C sky130_fd_sc_hd__nor2_1
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09914_ _09922_/A _09914_/B _09914_/C vssd1 vssd1 vccd1 vccd1 _09915_/A sky130_fd_sc_hd__and3_1
XFILLER_86_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09845_ _09845_/A vssd1 vssd1 vccd1 vccd1 _15433_/D sky130_fd_sc_hd__clkbuf_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09776_ _10065_/A vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08727_ _08724_/B _08724_/C _08726_/X vssd1 vssd1 vccd1 vccd1 _08728_/C sky130_fd_sc_hd__o21ai_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08658_ _15251_/Q _08657_/C _08590_/X vssd1 vssd1 vccd1 vccd1 _08659_/B sky130_fd_sc_hd__a21oi_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ state1[7] state1[6] state1[5] _07608_/X vssd1 vssd1 vccd1 vccd1 _15197_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _10969_/A vssd1 vssd1 vccd1 vccd1 _13078_/B sky130_fd_sc_hd__buf_2
X_10620_ _10627_/A _10618_/Y _10619_/Y _10615_/C vssd1 vssd1 vccd1 vccd1 _10622_/B
+ sky130_fd_sc_hd__o211a_1
X_10551_ _10549_/Y _10544_/C _10546_/X _10547_/Y vssd1 vssd1 vccd1 vccd1 _10552_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10482_ _10503_/A _10482_/B _10482_/C vssd1 vssd1 vccd1 vccd1 _10483_/A sky130_fd_sc_hd__and3_1
XFILLER_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13270_ _15976_/Q _13276_/C _13269_/X vssd1 vssd1 vccd1 vccd1 _13272_/C sky130_fd_sc_hd__a21o_1
X_12221_ _15806_/Q _12391_/B _12228_/C vssd1 vssd1 vccd1 vccd1 _12221_/X sky130_fd_sc_hd__and3_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ _12150_/X _12151_/Y _12147_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12154_/B
+ sky130_fd_sc_hd__o211ai_1
X_11103_ _11136_/C vssd1 vssd1 vccd1 vccd1 _11143_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12083_ _15784_/Q _12309_/B _12092_/C vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__and3_1
XFILLER_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11034_ _11612_/A vssd1 vssd1 vccd1 vccd1 _11267_/A sky130_fd_sc_hd__clkbuf_2
X_15911_ _15196_/Q _15911_/D vssd1 vssd1 vccd1 vccd1 _15911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15842_ _15907_/CLK _15842_/D vssd1 vssd1 vccd1 vccd1 _15842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15773_ _15890_/CLK _15773_/D vssd1 vssd1 vccd1 vccd1 _15773_/Q sky130_fd_sc_hd__dfxtp_1
X_12985_ _13004_/C vssd1 vssd1 vccd1 vccd1 _13016_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14724_ _14722_/A _14722_/B _14723_/X vssd1 vssd1 vccd1 vccd1 _16255_/D sky130_fd_sc_hd__a21oi_1
X_11936_ _15761_/Q _12107_/B _11943_/C vssd1 vssd1 vccd1 vccd1 _11936_/X sky130_fd_sc_hd__and3_1
XFILLER_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14655_ _07701_/X _14652_/A _07690_/X vssd1 vssd1 vccd1 vccd1 _14656_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ _11883_/A _11867_/B _11867_/C vssd1 vssd1 vccd1 vccd1 _11868_/A sky130_fd_sc_hd__and3_1
X_13606_ _16034_/Q _13605_/C _13452_/X vssd1 vssd1 vccd1 vccd1 _13607_/B sky130_fd_sc_hd__a21oi_1
X_10818_ _10931_/A _10818_/B _10822_/A vssd1 vssd1 vccd1 vccd1 _15585_/D sky130_fd_sc_hd__nor3_1
X_14586_ _14979_/A vssd1 vssd1 vccd1 vccd1 _14748_/A sky130_fd_sc_hd__buf_2
X_11798_ _12654_/A vssd1 vssd1 vccd1 vccd1 _11798_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16325_ _16327_/CLK _16325_/D vssd1 vssd1 vccd1 vccd1 _16325_/Q sky130_fd_sc_hd__dfxtp_2
X_13537_ _13529_/B _13530_/C _13533_/X _13535_/Y vssd1 vssd1 vccd1 vccd1 _13538_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10749_ _10978_/A vssd1 vssd1 vccd1 vccd1 _10789_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16256_ _16268_/CLK _16256_/D vssd1 vssd1 vccd1 vccd1 _16256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13468_ _16025_/Q _16024_/Q _16023_/Q _13467_/X vssd1 vssd1 vccd1 vccd1 _16008_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15207_ _16353_/CLK _15207_/D vssd1 vssd1 vccd1 vccd1 _15207_/Q sky130_fd_sc_hd__dfxtp_1
X_12419_ _15844_/Q _15843_/Q _15842_/Q _12418_/X vssd1 vssd1 vccd1 vccd1 _15836_/D
+ sky130_fd_sc_hd__o31a_1
X_16187_ _16187_/CLK _16187_/D vssd1 vssd1 vccd1 vccd1 _16187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13399_ _13476_/A _13399_/B _13404_/B vssd1 vssd1 vccd1 vccd1 _15995_/D sky130_fd_sc_hd__nor3_1
X_15138_ _16357_/Q _15142_/C _14988_/X vssd1 vssd1 vccd1 vccd1 _15138_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15069_ _15075_/A _15068_/Y _15064_/B _15065_/C vssd1 vssd1 vccd1 vccd1 _15071_/B
+ sky130_fd_sc_hd__o211a_1
X_07960_ _07960_/A vssd1 vssd1 vccd1 vccd1 _15061_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_4_clk _15584_/CLK vssd1 vssd1 vccd1 vccd1 _15230_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07891_ _07891_/A _07891_/B vssd1 vssd1 vccd1 vccd1 _07892_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09630_ _11128_/A vssd1 vssd1 vccd1 vccd1 _10785_/A sky130_fd_sc_hd__buf_4
XFILLER_56_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09561_ _09575_/A _09561_/B _09561_/C vssd1 vssd1 vccd1 vccd1 _09562_/A sky130_fd_sc_hd__and3_1
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08512_ _15231_/Q _11080_/A _08522_/C vssd1 vssd1 vccd1 vccd1 _08512_/X sky130_fd_sc_hd__and3_1
XFILLER_82_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09492_ _09493_/B _09493_/C _09493_/A vssd1 vssd1 vccd1 vccd1 _09494_/B sky130_fd_sc_hd__a21o_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08443_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08446_/A sky130_fd_sc_hd__nand2_1
X_08374_ _08331_/Y _08333_/X _08373_/Y vssd1 vssd1 vccd1 vccd1 _08375_/B sky130_fd_sc_hd__o21a_1
XFILLER_149_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09828_ _09865_/A _09828_/B _09828_/C vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__and3_1
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09759_ _09759_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09764_/C sky130_fd_sc_hd__nor2_1
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12804_/A _12770_/B _12774_/A vssd1 vssd1 vccd1 vccd1 _15891_/D sky130_fd_sc_hd__nor3_1
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11721_ _11727_/B _11721_/B vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__or2_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _16195_/Q _14440_/B _14447_/C vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__and3_1
X_11652_ _11650_/Y _11646_/C _11648_/X _11649_/Y vssd1 vssd1 vccd1 vccd1 _11653_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10603_ _15553_/Q _10604_/C _10373_/X vssd1 vssd1 vccd1 vccd1 _10603_/Y sky130_fd_sc_hd__a21oi_1
X_14371_ _14325_/X _14366_/B _14326_/X vssd1 vssd1 vccd1 vccd1 _14374_/A sky130_fd_sc_hd__a21oi_1
X_11583_ _15706_/Q _11811_/B _11585_/C vssd1 vssd1 vccd1 vccd1 _11583_/X sky130_fd_sc_hd__and3_1
X_16110_ _16129_/CLK _16110_/D vssd1 vssd1 vccd1 vccd1 _16110_/Q sky130_fd_sc_hd__dfxtp_2
X_13322_ _15985_/Q _13327_/C _13269_/X vssd1 vssd1 vccd1 vccd1 _13324_/C sky130_fd_sc_hd__a21o_1
X_10534_ _15542_/Q _10590_/B _10540_/C vssd1 vssd1 vccd1 vccd1 _10537_/B sky130_fd_sc_hd__nand3_1
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16041_ _16052_/CLK _16041_/D vssd1 vssd1 vccd1 vccd1 _16041_/Q sky130_fd_sc_hd__dfxtp_1
X_10465_ _10463_/B _10463_/C _10464_/X vssd1 vssd1 vccd1 vccd1 _10466_/C sky130_fd_sc_hd__o21ai_1
XFILLER_108_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13253_ _13457_/A _13255_/C vssd1 vssd1 vccd1 vccd1 _13253_/X sky130_fd_sc_hd__or2_1
XFILLER_108_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12204_ _12204_/A _12204_/B _12204_/C vssd1 vssd1 vccd1 vccd1 _12205_/C sky130_fd_sc_hd__nand3_1
X_10396_ _15520_/Q _10395_/C _10333_/X vssd1 vssd1 vccd1 vccd1 _10397_/B sky130_fd_sc_hd__a21oi_1
X_13184_ _13223_/A _13184_/B _13184_/C vssd1 vssd1 vccd1 vccd1 _13185_/A sky130_fd_sc_hd__and3_1
XFILLER_123_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12135_ _15797_/Q _15799_/Q _15798_/Q _12134_/X vssd1 vssd1 vccd1 vccd1 _15791_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_145_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12066_ _12066_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12067_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ _11014_/X _11015_/Y _11016_/Y _11011_/C vssd1 vssd1 vccd1 vccd1 _11019_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_65_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15825_ _15907_/CLK _15825_/D vssd1 vssd1 vccd1 vccd1 _15825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15756_ _15794_/CLK _15756_/D vssd1 vssd1 vccd1 vccd1 _15756_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ _15925_/Q _13078_/B _12968_/C vssd1 vssd1 vccd1 vccd1 _12977_/B sky130_fd_sc_hd__and3_1
XFILLER_33_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14707_ hold9/A _14706_/C _15165_/B vssd1 vssd1 vccd1 vccd1 _14709_/C sky130_fd_sc_hd__a21o_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11919_ _11919_/A _11919_/B _11919_/C vssd1 vssd1 vccd1 vccd1 _11920_/C sky130_fd_sc_hd__nand3_1
X_15687_ _15763_/CLK _15687_/D vssd1 vssd1 vccd1 vccd1 _15687_/Q sky130_fd_sc_hd__dfxtp_1
X_12899_ _12906_/A _12899_/B _12899_/C vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__and3_1
XFILLER_61_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14638_ _14716_/A _14638_/B _14642_/B vssd1 vssd1 vccd1 vccd1 _16236_/D sky130_fd_sc_hd__nor3_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14569_ _14565_/Y _14568_/X _14528_/X vssd1 vssd1 vccd1 vccd1 _14569_/Y sky130_fd_sc_hd__a21oi_1
X_16308_ _16312_/CLK _16308_/D vssd1 vssd1 vccd1 vccd1 _16308_/Q sky130_fd_sc_hd__dfxtp_2
X_08090_ _10058_/A _07751_/B _07750_/B vssd1 vssd1 vccd1 vccd1 _08096_/A sky130_fd_sc_hd__o21a_1
XFILLER_109_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16239_ _16268_/CLK _16239_/D vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _08999_/A _08992_/B _08992_/C vssd1 vssd1 vccd1 vccd1 _08993_/A sky130_fd_sc_hd__and3_1
XFILLER_102_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07943_ _08163_/A _07943_/B vssd1 vssd1 vccd1 vccd1 _08420_/C sky130_fd_sc_hd__or2_2
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07874_ _14584_/C _07874_/B vssd1 vssd1 vccd1 vccd1 _07991_/A sky130_fd_sc_hd__xnor2_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09613_ _09635_/A _09613_/B _09613_/C vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__and3_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09544_ _09557_/C vssd1 vssd1 vccd1 vccd1 _09565_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09475_ _10341_/A vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08426_ _08421_/C _08424_/Y _08425_/Y vssd1 vssd1 vccd1 vccd1 _15216_/D sky130_fd_sc_hd__o21a_1
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08357_ _08388_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__nor2_1
XFILLER_149_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08288_ _08198_/A _08198_/B _08287_/Y vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__a21o_1
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10250_ _10244_/B _10245_/C _10247_/X _10248_/Y vssd1 vssd1 vccd1 vccd1 _10251_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _16094_/Q _13945_/C _14587_/B vssd1 vssd1 vccd1 vccd1 _13942_/C sky130_fd_sc_hd__a21o_1
XFILLER_93_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13871_ _13885_/C vssd1 vssd1 vccd1 vccd1 _13903_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15610_ _15194_/Q _15610_/D vssd1 vssd1 vccd1 vccd1 _15610_/Q sky130_fd_sc_hd__dfxtp_1
X_12822_ _12854_/C vssd1 vssd1 vccd1 vccd1 _12861_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15541_ _15655_/CLK _15541_/D vssd1 vssd1 vccd1 vccd1 _15541_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _12919_/A _12757_/C vssd1 vssd1 vccd1 vccd1 _12753_/X sky130_fd_sc_hd__or2_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11704_ _12277_/A vssd1 vssd1 vccd1 vccd1 _11938_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _15483_/CLK _15472_/D vssd1 vssd1 vccd1 vccd1 _15472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _15879_/Q _12798_/B _12684_/C vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__and3_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14426_/C vssd1 vssd1 vccd1 vccd1 _14435_/C sky130_fd_sc_hd__clkbuf_1
X_11635_ _15714_/Q _11863_/B _11635_/C vssd1 vssd1 vccd1 vccd1 _11635_/X sky130_fd_sc_hd__and3_1
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14354_ _14353_/X _14352_/Y _14309_/X vssd1 vssd1 vccd1 vccd1 _14354_/Y sky130_fd_sc_hd__a21oi_1
X_11566_ _15703_/Q _11605_/C _11336_/X vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13305_ _14653_/A vssd1 vssd1 vccd1 vccd1 _13305_/X sky130_fd_sc_hd__clkbuf_2
X_10517_ _10629_/A _10520_/C vssd1 vssd1 vccd1 vccd1 _10517_/X sky130_fd_sc_hd__or2_1
XFILLER_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14285_ _14289_/C vssd1 vssd1 vccd1 vccd1 _14299_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_143_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11497_ _11727_/A _11497_/B _11497_/C vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__or3_1
XFILLER_109_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16024_ _16040_/CLK _16024_/D vssd1 vssd1 vccd1 vccd1 _16024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ _13234_/Y _13230_/C _13232_/X _13233_/Y vssd1 vssd1 vccd1 vccd1 _13237_/C
+ sky130_fd_sc_hd__a211o_1
X_10448_ _10736_/A vssd1 vssd1 vccd1 vccd1 _10681_/B sky130_fd_sc_hd__buf_2
XFILLER_124_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _15958_/Q _13172_/C _14250_/A vssd1 vssd1 vccd1 vccd1 _13169_/C sky130_fd_sc_hd__a21o_1
X_10379_ _10379_/A vssd1 vssd1 vccd1 vccd1 _15516_/D sky130_fd_sc_hd__clkbuf_1
X_12118_ _12124_/A _12116_/Y _12117_/Y _12112_/C vssd1 vssd1 vccd1 vccd1 _12120_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13098_ _13218_/A _13098_/B _13105_/A vssd1 vssd1 vccd1 vccd1 _15946_/D sky130_fd_sc_hd__nor3_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12049_ _15779_/Q _12055_/C _12048_/X vssd1 vssd1 vccd1 vccd1 _12049_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15808_ _07603_/A _15808_/D vssd1 vssd1 vccd1 vccd1 _15808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15739_ _15794_/CLK _15739_/D vssd1 vssd1 vccd1 vccd1 _15739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ _15344_/Q _09297_/C _09029_/X vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__a21oi_1
X_08211_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08211_/Y sky130_fd_sc_hd__xnor2_1
X_09191_ _09190_/B _09190_/C _09019_/X vssd1 vssd1 vccd1 vccd1 _09192_/C sky130_fd_sc_hd__o21ai_1
XFILLER_147_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08142_ _08256_/A _08256_/B vssd1 vssd1 vccd1 vccd1 _08143_/B sky130_fd_sc_hd__xor2_4
XFILLER_146_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08073_ _11213_/A _11332_/A _08072_/Y vssd1 vssd1 vccd1 vccd1 _08226_/B sky130_fd_sc_hd__o21ai_4
XFILLER_119_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08975_ _08976_/B _08976_/C _08976_/A vssd1 vssd1 vccd1 vccd1 _08977_/B sky130_fd_sc_hd__a21o_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_07926_ _15746_/Q _16341_/Q vssd1 vssd1 vccd1 vccd1 _07928_/A sky130_fd_sc_hd__or2_1
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07857_ _13729_/C _07857_/B vssd1 vssd1 vccd1 vccd1 _07859_/B sky130_fd_sc_hd__xnor2_4
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07788_ _15512_/Q vssd1 vssd1 vccd1 vccd1 _10347_/A sky130_fd_sc_hd__inv_2
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09527_ _09643_/A _09527_/B _09531_/B vssd1 vssd1 vccd1 vccd1 _15383_/D sky130_fd_sc_hd__nor3_1
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09458_ _09458_/A _09458_/B _09458_/C vssd1 vssd1 vccd1 vccd1 _09459_/A sky130_fd_sc_hd__and3_1
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08409_ _08415_/A _08468_/A vssd1 vssd1 vccd1 vccd1 _08411_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09389_ _13532_/A vssd1 vssd1 vccd1 vccd1 _10548_/A sky130_fd_sc_hd__buf_2
X_11420_ _11420_/A _11420_/B _11420_/C vssd1 vssd1 vccd1 vccd1 _11421_/A sky130_fd_sc_hd__and3_1
XFILLER_137_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ _11365_/A _11351_/B _11351_/C vssd1 vssd1 vccd1 vccd1 _11352_/A sky130_fd_sc_hd__and3_1
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10302_ _10323_/A _10302_/B _10302_/C vssd1 vssd1 vccd1 vccd1 _10303_/A sky130_fd_sc_hd__and3_1
X_14070_ _16119_/Q _14099_/C _14069_/X vssd1 vssd1 vccd1 vccd1 _14072_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11282_ _11569_/A vssd1 vssd1 vccd1 vccd1 _11510_/B sky130_fd_sc_hd__buf_2
XFILLER_118_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13021_ _13077_/A _13021_/B _13025_/B vssd1 vssd1 vccd1 vccd1 _15932_/D sky130_fd_sc_hd__nor3_1
X_10233_ _10388_/A vssd1 vssd1 vccd1 vccd1 _10353_/A sky130_fd_sc_hd__buf_2
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10164_ _10171_/B _10164_/B vssd1 vssd1 vccd1 vccd1 _10166_/A sky130_fd_sc_hd__or2_1
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10095_ _10092_/X _10093_/Y _10094_/Y _10088_/C vssd1 vssd1 vccd1 vccd1 _10097_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14972_ _14814_/X _14969_/A _14971_/Y vssd1 vssd1 vccd1 vccd1 _16313_/D sky130_fd_sc_hd__o21a_1
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13923_ _13921_/X _13917_/B _13922_/X vssd1 vssd1 vccd1 vccd1 _13923_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13854_ _16079_/Q _13853_/C _13708_/X vssd1 vssd1 vccd1 vccd1 _13855_/B sky130_fd_sc_hd__a21oi_1
XFILLER_142_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ _15898_/Q _12861_/B _12805_/C vssd1 vssd1 vccd1 vccd1 _12813_/B sky130_fd_sc_hd__and3_1
X_13785_ _16067_/Q _14080_/B _13785_/C vssd1 vssd1 vccd1 vccd1 _13785_/X sky130_fd_sc_hd__and3_1
X_10997_ _11019_/A _10997_/B _10997_/C vssd1 vssd1 vccd1 vccd1 _10998_/A sky130_fd_sc_hd__and3_1
X_15524_ _15655_/CLK _15524_/D vssd1 vssd1 vccd1 vccd1 _15524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _15887_/Q _12742_/C _12616_/X vssd1 vssd1 vccd1 vccd1 _12736_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ _15484_/CLK _15455_/D vssd1 vssd1 vccd1 vccd1 _15455_/Q sky130_fd_sc_hd__dfxtp_1
X_12667_ _15877_/Q _12667_/B _12670_/C vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__and3_1
X_14406_ _14401_/Y _14405_/X _14316_/X vssd1 vssd1 vccd1 vccd1 _14406_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11618_ _11618_/A vssd1 vssd1 vccd1 vccd1 _15709_/D sky130_fd_sc_hd__clkbuf_1
X_15386_ _15395_/CLK _15386_/D vssd1 vssd1 vccd1 vccd1 _15386_/Q sky130_fd_sc_hd__dfxtp_1
X_12598_ _12598_/A _12598_/B _12598_/C vssd1 vssd1 vccd1 vccd1 _12599_/C sky130_fd_sc_hd__nand3_1
X_14337_ _16174_/Q _14337_/B _14337_/C vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__and3_1
X_11549_ _11556_/B _11549_/B vssd1 vssd1 vccd1 vccd1 _11552_/A sky130_fd_sc_hd__or2_1
XFILLER_116_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14268_ _14265_/B _14264_/Y _14265_/A vssd1 vssd1 vccd1 vccd1 _14268_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_109_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16007_ _16007_/CLK _16007_/D vssd1 vssd1 vccd1 vccd1 _16007_/Q sky130_fd_sc_hd__dfxtp_1
X_13219_ _15967_/Q _13374_/B _13226_/C vssd1 vssd1 vccd1 vccd1 _13222_/B sky130_fd_sc_hd__nand3_1
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14199_ _14058_/X _14193_/B _14059_/X vssd1 vssd1 vccd1 vccd1 _14201_/A sky130_fd_sc_hd__a21oi_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08760_ _13640_/A vssd1 vssd1 vccd1 vccd1 _13693_/A sky130_fd_sc_hd__buf_6
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ _13930_/A vssd1 vssd1 vccd1 vccd1 _15181_/A sky130_fd_sc_hd__clkbuf_2
X_08691_ _08691_/A vssd1 vssd1 vccd1 vccd1 _15255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07642_ _12661_/A vssd1 vssd1 vccd1 vccd1 _12609_/A sky130_fd_sc_hd__buf_4
XFILLER_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09312_ _15342_/Q vssd1 vssd1 vccd1 vccd1 _09326_/C sky130_fd_sc_hd__inv_2
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09243_ _15341_/Q _09242_/C _09180_/X vssd1 vssd1 vccd1 vccd1 _09244_/B sky130_fd_sc_hd__a21oi_1
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09174_ _15331_/Q _09179_/C _09118_/X vssd1 vssd1 vccd1 vccd1 _09174_/Y sky130_fd_sc_hd__a21oi_1
X_08125_ _15243_/Q _08125_/B vssd1 vssd1 vccd1 vccd1 _08125_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08056_ _15737_/Q _08056_/B vssd1 vssd1 vccd1 vccd1 _08056_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08958_ _09185_/A _08961_/C vssd1 vssd1 vccd1 vccd1 _08958_/X sky130_fd_sc_hd__or2_1
XFILLER_69_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07909_ _07909_/A _07909_/B vssd1 vssd1 vccd1 vccd1 _07957_/B sky130_fd_sc_hd__xor2_4
X_08889_ _15287_/Q _08886_/C _08888_/X vssd1 vssd1 vccd1 vccd1 _08890_/B sky130_fd_sc_hd__a21oi_1
XFILLER_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10920_ _11151_/A _10920_/B _10920_/C vssd1 vssd1 vccd1 vccd1 _10922_/B sky130_fd_sc_hd__or3_1
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _10858_/A _10849_/Y _10850_/Y _10845_/C vssd1 vssd1 vccd1 vccd1 _10853_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _13575_/C vssd1 vssd1 vccd1 vccd1 _13583_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10782_ _10782_/A vssd1 vssd1 vccd1 vccd1 _15579_/D sky130_fd_sc_hd__clkbuf_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12527_/B _12521_/B vssd1 vssd1 vccd1 vccd1 _12523_/A sky130_fd_sc_hd__or2_1
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15351_/CLK _15240_/D vssd1 vssd1 vccd1 vccd1 _15240_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _12449_/X _12450_/Y _12451_/Y _12446_/C vssd1 vssd1 vccd1 vccd1 _12454_/B
+ sky130_fd_sc_hd__o211ai_1
X_11403_ _11401_/X _11402_/Y _11398_/B _11399_/C vssd1 vssd1 vccd1 vccd1 _11405_/B
+ sky130_fd_sc_hd__o211ai_1
X_15171_ _16366_/Q _15171_/B _15176_/C vssd1 vssd1 vccd1 vccd1 _15179_/A sky130_fd_sc_hd__and3_1
X_12383_ _15832_/Q _12383_/B _12386_/C vssd1 vssd1 vccd1 vccd1 _12383_/X sky130_fd_sc_hd__and3_1
X_14122_ _14122_/A _14122_/B _14122_/C vssd1 vssd1 vccd1 vccd1 _14123_/C sky130_fd_sc_hd__nand3_1
X_11334_ _11355_/C vssd1 vssd1 vccd1 vccd1 _11367_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14053_ _15186_/A _14053_/B vssd1 vssd1 vccd1 vccd1 _14054_/B sky130_fd_sc_hd__and2_1
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ _11493_/A _11268_/C vssd1 vssd1 vccd1 vccd1 _11265_/X sky130_fd_sc_hd__or2_1
XFILLER_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13004_ _15930_/Q _14031_/A _13004_/C vssd1 vssd1 vccd1 vccd1 _13004_/Y sky130_fd_sc_hd__nand3_1
X_10216_ _15491_/Q _10391_/B _10220_/C vssd1 vssd1 vccd1 vccd1 _10216_/Y sky130_fd_sc_hd__nand3_1
X_11196_ _11220_/A _11196_/B _11202_/B vssd1 vssd1 vccd1 vccd1 _15644_/D sky130_fd_sc_hd__nor3_1
XFILLER_95_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _10147_/A vssd1 vssd1 vccd1 vccd1 _15480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14955_ _14955_/A _14955_/B vssd1 vssd1 vccd1 vccd1 _14957_/A sky130_fd_sc_hd__or2_1
X_10078_ _10071_/B _10072_/C _10074_/X _10076_/Y vssd1 vssd1 vccd1 vccd1 _10079_/C
+ sky130_fd_sc_hd__a211o_1
X_13906_ _13903_/X _13906_/B vssd1 vssd1 vccd1 vccd1 _13906_/X sky130_fd_sc_hd__and2b_1
X_14886_ _14802_/X _14877_/A _14881_/B _14885_/Y vssd1 vssd1 vccd1 vccd1 _16292_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13837_ _13837_/A vssd1 vssd1 vccd1 vccd1 _16074_/D sky130_fd_sc_hd__clkbuf_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13768_ _13789_/A _13768_/B _13768_/C vssd1 vssd1 vccd1 vccd1 _13769_/A sky130_fd_sc_hd__and3_1
XFILLER_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15507_ _15224_/Q _15507_/D vssd1 vssd1 vccd1 vccd1 _15507_/Q sky130_fd_sc_hd__dfxtp_1
X_12719_ _12719_/A vssd1 vssd1 vccd1 vccd1 _15883_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_13699_ _13699_/A vssd1 vssd1 vccd1 vccd1 _16048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15438_ _15484_/CLK _15438_/D vssd1 vssd1 vccd1 vccd1 _15438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _15484_/CLK _15369_/D vssd1 vssd1 vccd1 vccd1 _15369_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09930_ _09930_/A _09930_/B _09934_/B vssd1 vssd1 vccd1 vccd1 _15446_/D sky130_fd_sc_hd__nor3_1
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09861_ _15437_/Q _09867_/C _09741_/X vssd1 vssd1 vccd1 vccd1 _09861_/Y sky130_fd_sc_hd__a21oi_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _08808_/X _08809_/Y _08811_/Y _08806_/C vssd1 vssd1 vccd1 vccd1 _08814_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_100_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _10081_/A vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08765_/A _08743_/B _08743_/C vssd1 vssd1 vccd1 vccd1 _08744_/A sky130_fd_sc_hd__and3_1
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08674_ _08694_/C vssd1 vssd1 vccd1 vccd1 _08706_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _15202_/Q _13316_/A _07633_/C vssd1 vssd1 vccd1 vccd1 _07638_/A sky130_fd_sc_hd__and3_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09226_ _09226_/A vssd1 vssd1 vccd1 vccd1 _15337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09157_ _09157_/A vssd1 vssd1 vccd1 vccd1 _15327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08108_ _07752_/A _07752_/B _08107_/X vssd1 vssd1 vccd1 vccd1 _08116_/A sky130_fd_sc_hd__o21a_1
X_09088_ _15317_/Q _09088_/B _09096_/C vssd1 vssd1 vccd1 vccd1 _09093_/A sky130_fd_sc_hd__and3_1
XFILLER_135_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08039_ _11156_/A _07848_/B _08038_/X vssd1 vssd1 vccd1 vccd1 _08201_/B sky130_fd_sc_hd__o21a_2
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11050_ _11085_/A _11050_/B _11054_/A vssd1 vssd1 vccd1 vccd1 _15621_/D sky130_fd_sc_hd__nor3_1
XFILLER_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10001_ _15466_/Q _15465_/Q _15464_/Q _09831_/X vssd1 vssd1 vccd1 vccd1 _15458_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14740_ _16265_/Q _14755_/C _14702_/X vssd1 vssd1 vccd1 vccd1 _14742_/B sky130_fd_sc_hd__a21oi_1
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11952_ _11958_/B _11952_/B vssd1 vssd1 vccd1 vccd1 _11954_/A sky130_fd_sc_hd__or2_1
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10903_ _10903_/A vssd1 vssd1 vccd1 vccd1 _15598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14671_ _14869_/A vssd1 vssd1 vccd1 vccd1 _14833_/B sky130_fd_sc_hd__buf_2
X_11883_ _11883_/A _11883_/B _11883_/C vssd1 vssd1 vccd1 vccd1 _11884_/A sky130_fd_sc_hd__and3_1
X_13622_ _13626_/C vssd1 vssd1 vccd1 vccd1 _13634_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10834_ _12041_/A vssd1 vssd1 vccd1 vccd1 _11121_/B sky130_fd_sc_hd__buf_2
XFILLER_32_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater13 _15195_/Q vssd1 vssd1 vccd1 vccd1 _15794_/CLK sky130_fd_sc_hd__buf_12
X_16341_ _16352_/CLK _16341_/D vssd1 vssd1 vccd1 vccd1 _16341_/Q sky130_fd_sc_hd__dfxtp_1
X_13553_ _13604_/A _13553_/B _13557_/B vssd1 vssd1 vccd1 vccd1 _16022_/D sky130_fd_sc_hd__nor3_1
X_10765_ _15578_/Q _10770_/C _10648_/X vssd1 vssd1 vccd1 vccd1 _10767_/C sky130_fd_sc_hd__a21o_1
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ _12504_/A vssd1 vssd1 vccd1 vccd1 _15849_/D sky130_fd_sc_hd__clkbuf_1
X_16272_ _16273_/CLK _16272_/D vssd1 vssd1 vccd1 vccd1 _16272_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13484_ _16013_/Q _13484_/B _13484_/C vssd1 vssd1 vccd1 vccd1 _13484_/X sky130_fd_sc_hd__and3_1
X_10696_ _10732_/A _10696_/B _10696_/C vssd1 vssd1 vccd1 vccd1 _10697_/A sky130_fd_sc_hd__and3_1
X_15223_ _15260_/CLK _15223_/D vssd1 vssd1 vccd1 vccd1 _15223_/Q sky130_fd_sc_hd__dfxtp_1
X_12435_ _15840_/Q _12443_/C _12377_/X vssd1 vssd1 vccd1 vccd1 _12435_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15154_ _15154_/A _15154_/B vssd1 vssd1 vccd1 vccd1 _16356_/D sky130_fd_sc_hd__nor2_1
XFILLER_126_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12366_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12593_/B sky130_fd_sc_hd__buf_2
X_14105_ _14103_/A _14103_/B _14104_/X vssd1 vssd1 vccd1 vccd1 _16122_/D sky130_fd_sc_hd__a21oi_1
X_11317_ _15664_/Q _11431_/B _11317_/C vssd1 vssd1 vccd1 vccd1 _11326_/B sky130_fd_sc_hd__and3_1
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15085_ _15189_/A _15189_/B _15085_/C vssd1 vssd1 vccd1 vccd1 _15088_/A sky130_fd_sc_hd__and3_1
XFILLER_126_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12297_ _12295_/A _12295_/B _12296_/X vssd1 vssd1 vccd1 vccd1 _15816_/D sky130_fd_sc_hd__a21oi_1
XFILLER_141_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14036_ _14028_/B _14029_/C _14040_/A _14034_/Y vssd1 vssd1 vccd1 vccd1 _14040_/B
+ sky130_fd_sc_hd__a211oi_1
X_11248_ _11246_/Y _11242_/C _11244_/X _11245_/Y vssd1 vssd1 vccd1 vccd1 _11249_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ _11175_/X _11176_/Y _11178_/Y _11173_/C vssd1 vssd1 vccd1 vccd1 _11181_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_121_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15987_ _16052_/CLK _15987_/D vssd1 vssd1 vccd1 vccd1 _15987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14938_ _16310_/Q _14953_/C _14901_/X vssd1 vssd1 vccd1 vccd1 _14940_/B sky130_fd_sc_hd__a21oi_1
X_14869_ _14869_/A vssd1 vssd1 vccd1 vccd1 _15031_/B sky130_fd_sc_hd__buf_2
XFILLER_51_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08390_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08393_/A sky130_fd_sc_hd__xor2_4
XFILLER_16_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09011_ _09011_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _09012_/B sky130_fd_sc_hd__nor2_1
XFILLER_117_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09913_ _09911_/Y _09907_/C _09909_/X _09910_/Y vssd1 vssd1 vccd1 vccd1 _09914_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _09865_/A _09844_/B _09844_/C vssd1 vssd1 vccd1 vccd1 _09845_/A sky130_fd_sc_hd__and3_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _09775_/A _09775_/B _09781_/A vssd1 vssd1 vccd1 vccd1 _15423_/D sky130_fd_sc_hd__nor3_1
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08726_ _14372_/A vssd1 vssd1 vccd1 vccd1 _08726_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _15251_/Q _08775_/B _08657_/C vssd1 vssd1 vccd1 vccd1 _08667_/B sky130_fd_sc_hd__and3_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _09541_/A vssd1 vssd1 vccd1 vccd1 _07608_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08588_ _15242_/Q _08775_/B _08588_/C vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__and3_1
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10550_ _10546_/X _10547_/Y _10549_/Y _10544_/C vssd1 vssd1 vccd1 vccd1 _10552_/B
+ sky130_fd_sc_hd__o211ai_1
X_09209_ _09233_/A _09209_/B _09209_/C vssd1 vssd1 vccd1 vccd1 _09210_/A sky130_fd_sc_hd__and3_1
X_10481_ _10481_/A _10481_/B _10481_/C vssd1 vssd1 vccd1 vccd1 _10482_/C sky130_fd_sc_hd__nand3_1
XFILLER_108_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ _12220_/A vssd1 vssd1 vccd1 vccd1 _15804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ _15795_/Q _12159_/C _12093_/X vssd1 vssd1 vccd1 vccd1 _12151_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11102_ _11121_/C vssd1 vssd1 vccd1 vccd1 _11136_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12082_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12309_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_1_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11033_ _11031_/A _11031_/B _11032_/X vssd1 vssd1 vccd1 vccd1 _15618_/D sky130_fd_sc_hd__a21oi_1
X_15910_ _15196_/Q _15910_/D vssd1 vssd1 vccd1 vccd1 _15910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15841_ _15907_/CLK _15841_/D vssd1 vssd1 vccd1 vccd1 _15841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15772_ _15195_/Q _15772_/D vssd1 vssd1 vccd1 vccd1 _15772_/Q sky130_fd_sc_hd__dfxtp_1
X_12984_ _12996_/C vssd1 vssd1 vccd1 vccd1 _13004_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11935_ _11935_/A vssd1 vssd1 vccd1 vccd1 _15759_/D sky130_fd_sc_hd__clkbuf_1
X_14723_ _14843_/A _14723_/B vssd1 vssd1 vccd1 vccd1 _14723_/X sky130_fd_sc_hd__or2_1
XFILLER_33_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14654_ _14964_/A _14811_/B _14654_/C vssd1 vssd1 vccd1 vccd1 _14656_/A sky130_fd_sc_hd__and3_1
X_11866_ _11860_/B _11861_/C _11863_/X _11864_/Y vssd1 vssd1 vccd1 vccd1 _11867_/C
+ sky130_fd_sc_hd__a211o_1
X_13605_ _16034_/Q _13605_/B _13605_/C vssd1 vssd1 vccd1 vccd1 _13613_/B sky130_fd_sc_hd__and3_1
X_10817_ _15586_/Q _10817_/B _10825_/C vssd1 vssd1 vccd1 vccd1 _10822_/A sky130_fd_sc_hd__and3_1
X_14585_ _14626_/A _14585_/B _14590_/A vssd1 vssd1 vccd1 vccd1 _16225_/D sky130_fd_sc_hd__nor3_1
X_11797_ _15740_/Q _11797_/B _11804_/C vssd1 vssd1 vccd1 vccd1 _11801_/B sky130_fd_sc_hd__nand3_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13536_ _13533_/X _13535_/Y _13529_/B _13530_/C vssd1 vssd1 vccd1 vccd1 _13538_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16324_ _16327_/CLK _16324_/D vssd1 vssd1 vccd1 vccd1 _16324_/Q sky130_fd_sc_hd__dfxtp_2
X_10748_ _11612_/A vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16255_ _16264_/CLK _16255_/D vssd1 vssd1 vccd1 vccd1 _16255_/Q sky130_fd_sc_hd__dfxtp_2
X_13467_ _13723_/A vssd1 vssd1 vccd1 vccd1 _13467_/X sky130_fd_sc_hd__clkbuf_2
X_10679_ _15564_/Q _10734_/B _10679_/C vssd1 vssd1 vccd1 vccd1 _10688_/A sky130_fd_sc_hd__and3_1
X_15206_ _16353_/CLK _15206_/D vssd1 vssd1 vccd1 vccd1 _15206_/Q sky130_fd_sc_hd__dfxtp_2
X_12418_ _12418_/A vssd1 vssd1 vccd1 vccd1 _12418_/X sky130_fd_sc_hd__buf_2
XFILLER_127_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16186_ _16187_/CLK _16186_/D vssd1 vssd1 vccd1 vccd1 _16186_/Q sky130_fd_sc_hd__dfxtp_1
X_13398_ _13396_/Y _13392_/C _13404_/A _13395_/Y vssd1 vssd1 vccd1 vccd1 _13404_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ _16357_/Q _15171_/B _15142_/C vssd1 vssd1 vccd1 vccd1 _15145_/A sky130_fd_sc_hd__and3_1
X_12349_ _12356_/B _12349_/B vssd1 vssd1 vccd1 vccd1 _12351_/A sky130_fd_sc_hd__or2_1
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15068_ _16339_/Q _15072_/C _14988_/X vssd1 vssd1 vccd1 vccd1 _15068_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14019_ _14022_/C vssd1 vssd1 vccd1 vccd1 _14032_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07890_ _15422_/Q _07890_/B vssd1 vssd1 vccd1 vccd1 _07891_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09560_ _09553_/B _09554_/C _09557_/X _09558_/Y vssd1 vssd1 vccd1 vccd1 _09561_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_83_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08511_ _10896_/A vssd1 vssd1 vccd1 vccd1 _11080_/A sky130_fd_sc_hd__buf_4
XFILLER_64_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09491_ _15380_/Q _09496_/C _09490_/X vssd1 vssd1 vccd1 vccd1 _09493_/C sky130_fd_sc_hd__a21o_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08442_ _08442_/A _08442_/B vssd1 vssd1 vccd1 vccd1 _08443_/B sky130_fd_sc_hd__or2_1
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08373_ _08373_/A _08444_/A vssd1 vssd1 vccd1 vccd1 _08373_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09827_ _09826_/B _09826_/C _09596_/X vssd1 vssd1 vccd1 vccd1 _09828_/C sky130_fd_sc_hd__o21ai_1
XFILLER_48_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09758_ _09758_/A _09758_/B vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__nor2_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ _13700_/A vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__buf_6
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _09687_/Y _09683_/C _09685_/X _09686_/Y vssd1 vssd1 vccd1 vccd1 _09690_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_64_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _15727_/Q _11719_/C _11488_/X vssd1 vssd1 vccd1 vccd1 _11721_/B sky130_fd_sc_hd__a21oi_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11651_ _11648_/X _11649_/Y _11650_/Y _11646_/C vssd1 vssd1 vccd1 vccd1 _11653_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10602_ _15553_/Q _10602_/B _10604_/C vssd1 vssd1 vccd1 vccd1 _10602_/X sky130_fd_sc_hd__and3_1
X_14370_ _14195_/X _14366_/B _14369_/Y vssd1 vssd1 vccd1 vccd1 _16177_/D sky130_fd_sc_hd__o21a_1
X_11582_ _11582_/A vssd1 vssd1 vccd1 vccd1 _11811_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13321_ _15985_/Q _13374_/B _13327_/C vssd1 vssd1 vccd1 vccd1 _13324_/B sky130_fd_sc_hd__nand3_1
X_10533_ _10645_/A _10533_/B _10537_/A vssd1 vssd1 vccd1 vccd1 _15540_/D sky130_fd_sc_hd__nor3_1
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16040_ _16040_/CLK _16040_/D vssd1 vssd1 vccd1 vccd1 _16040_/Q sky130_fd_sc_hd__dfxtp_1
X_13252_ _13252_/A _13252_/B vssd1 vssd1 vccd1 vccd1 _13255_/C sky130_fd_sc_hd__nor2_1
X_10464_ _10751_/A vssd1 vssd1 vccd1 vccd1 _10464_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ _12204_/B _12204_/C _12204_/A vssd1 vssd1 vccd1 vccd1 _12205_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13183_ _13181_/Y _13176_/C _13178_/X _13180_/Y vssd1 vssd1 vccd1 vccd1 _13184_/C
+ sky130_fd_sc_hd__a211o_1
X_10395_ _15520_/Q _10512_/B _10395_/C vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__and3_1
XFILLER_123_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _12418_/A vssd1 vssd1 vccd1 vccd1 _12134_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12065_ _12072_/B _12065_/B vssd1 vssd1 vccd1 vccd1 _12067_/A sky130_fd_sc_hd__or2_1
X_11016_ _15616_/Q _11073_/B _11021_/C vssd1 vssd1 vccd1 vccd1 _11016_/Y sky130_fd_sc_hd__nand3_1
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15824_ _15907_/CLK _15824_/D vssd1 vssd1 vccd1 vccd1 _15824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15755_ _15890_/CLK _15755_/D vssd1 vssd1 vccd1 vccd1 _15755_/Q sky130_fd_sc_hd__dfxtp_1
X_12967_ _13077_/A _12967_/B _12971_/B vssd1 vssd1 vccd1 vccd1 _15923_/D sky130_fd_sc_hd__nor3_1
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11918_ _11919_/B _11919_/C _11919_/A vssd1 vssd1 vccd1 vccd1 _11920_/B sky130_fd_sc_hd__a21o_1
X_14706_ hold9/A _14743_/B _14706_/C vssd1 vssd1 vccd1 vccd1 _14709_/B sky130_fd_sc_hd__nand3_1
X_15686_ _15763_/CLK _15686_/D vssd1 vssd1 vccd1 vccd1 _15686_/Q sky130_fd_sc_hd__dfxtp_1
X_12898_ _12896_/Y _12891_/C _12893_/X _12894_/Y vssd1 vssd1 vccd1 vccd1 _12899_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11849_ _15746_/Q vssd1 vssd1 vccd1 vccd1 _11863_/C sky130_fd_sc_hd__inv_2
X_14637_ _14630_/B _14631_/C _14642_/A _14635_/Y vssd1 vssd1 vccd1 vccd1 _14642_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _14566_/X _14568_/B vssd1 vssd1 vccd1 vccd1 _14568_/X sky130_fd_sc_hd__and2b_1
X_16307_ _16312_/CLK _16307_/D vssd1 vssd1 vccd1 vccd1 _16307_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13519_ _13523_/C vssd1 vssd1 vccd1 vccd1 _13533_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14499_ _14499_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _16205_/D sky130_fd_sc_hd__nor2_1
X_16238_ _16247_/CLK _16238_/D vssd1 vssd1 vccd1 vccd1 _16238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16169_ _16169_/CLK _16169_/D vssd1 vssd1 vccd1 vccd1 _16169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08991_ _08989_/Y _08985_/C _08987_/X _08988_/Y vssd1 vssd1 vccd1 vccd1 _08992_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_142_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07942_ _08622_/C _07942_/B vssd1 vssd1 vccd1 vccd1 _07943_/B sky130_fd_sc_hd__and2_1
XFILLER_102_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07873_ _07873_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07874_/B sky130_fd_sc_hd__nand2_2
XFILLER_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09612_ _09612_/A _09612_/B _09612_/C vssd1 vssd1 vccd1 vccd1 _09613_/C sky130_fd_sc_hd__nand3_1
XFILLER_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09543_ _09543_/A vssd1 vssd1 vccd1 vccd1 _09557_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09474_ _09536_/A vssd1 vssd1 vccd1 vccd1 _09519_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08425_ _08421_/C _08424_/Y _08168_/X vssd1 vssd1 vccd1 vccd1 _08425_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08356_ _08356_/A _08356_/B _08356_/C vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__and3_1
XFILLER_149_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08287_ _08287_/A _08287_/B vssd1 vssd1 vccd1 vccd1 _08287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10180_ _10214_/C vssd1 vssd1 vccd1 vccd1 _10220_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13870_ _13874_/C vssd1 vssd1 vccd1 vccd1 _13885_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _12840_/C vssd1 vssd1 vccd1 vccd1 _12854_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15540_ _15655_/CLK _15540_/D vssd1 vssd1 vccd1 vccd1 _15540_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _12752_/A _12752_/B vssd1 vssd1 vccd1 vccd1 _12757_/C sky130_fd_sc_hd__nor2_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _15725_/Q _11712_/C _11472_/X vssd1 vssd1 vccd1 vccd1 _11703_/Y sky130_fd_sc_hd__a21oi_1
X_15471_ _15483_/CLK _15471_/D vssd1 vssd1 vccd1 vccd1 _15471_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12683_ _13239_/A vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__buf_2
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _16205_/Q _16204_/Q _16203_/Q _14421_/X vssd1 vssd1 vccd1 vccd1 _16188_/D
+ sky130_fd_sc_hd__o31a_1
X_11634_ _11634_/A vssd1 vssd1 vccd1 vccd1 _11863_/B sky130_fd_sc_hd__clkbuf_2
X_16375__24 vssd1 vssd1 vccd1 vccd1 _16375__24/HI io_oeb[7] sky130_fd_sc_hd__conb_1
XFILLER_11_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14353_ _14353_/A _14353_/B vssd1 vssd1 vccd1 vccd1 _14353_/X sky130_fd_sc_hd__or2_1
XFILLER_11_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11565_ _11599_/C vssd1 vssd1 vccd1 vccd1 _11605_/C sky130_fd_sc_hd__clkbuf_2
X_13304_ _13408_/A _13304_/B _13304_/C vssd1 vssd1 vccd1 vccd1 _13307_/B sky130_fd_sc_hd__or3_1
X_10516_ _10516_/A _10516_/B vssd1 vssd1 vccd1 vccd1 _10520_/C sky130_fd_sc_hd__nor2_1
XFILLER_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14284_ _16178_/Q _16177_/Q _16176_/Q _14202_/X vssd1 vssd1 vccd1 vccd1 _16161_/D
+ sky130_fd_sc_hd__o31a_1
X_11496_ _11783_/A vssd1 vssd1 vccd1 vccd1 _11727_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13235_ _13232_/X _13233_/Y _13234_/Y _13230_/C vssd1 vssd1 vccd1 vccd1 _13237_/B
+ sky130_fd_sc_hd__o211ai_1
X_16023_ _16031_/CLK _16023_/D vssd1 vssd1 vccd1 vccd1 _16023_/Q sky130_fd_sc_hd__dfxtp_1
X_10447_ _15528_/Q _10453_/C _10269_/X vssd1 vssd1 vccd1 vccd1 _10447_/Y sky130_fd_sc_hd__a21oi_1
X_13166_ _15958_/Q _13374_/B _13172_/C vssd1 vssd1 vccd1 vccd1 _13169_/B sky130_fd_sc_hd__nand3_1
X_10378_ _10386_/A _10378_/B _10378_/C vssd1 vssd1 vccd1 vccd1 _10379_/A sky130_fd_sc_hd__and3_1
X_12117_ _15788_/Q _12174_/B _12121_/C vssd1 vssd1 vccd1 vccd1 _12117_/Y sky130_fd_sc_hd__nand3_1
XFILLER_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13097_ _15948_/Q _14379_/A _13097_/C vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__and3_1
X_12048_ _12048_/A vssd1 vssd1 vccd1 vccd1 _12048_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15807_ _07603_/A _15807_/D vssd1 vssd1 vccd1 vccd1 _15807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13999_ _13999_/A _13999_/B vssd1 vssd1 vccd1 vccd1 _13999_/X sky130_fd_sc_hd__or2_1
XFILLER_34_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15738_ _15794_/CLK _15738_/D vssd1 vssd1 vccd1 vccd1 _15738_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15669_ _15763_/CLK _15669_/D vssd1 vssd1 vccd1 vccd1 _15669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08210_ _08035_/A _08035_/B _08034_/A vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__a21oi_4
X_09190_ _09419_/A _09190_/B _09190_/C vssd1 vssd1 vccd1 vccd1 _09192_/B sky130_fd_sc_hd__or3_1
XFILLER_147_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08141_ _07786_/A _07786_/B _08140_/Y vssd1 vssd1 vccd1 vccd1 _08256_/B sky130_fd_sc_hd__o21a_2
XFILLER_146_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08072_ _15683_/Q _08072_/B vssd1 vssd1 vccd1 vccd1 _08072_/Y sky130_fd_sc_hd__nand2_1
XFILLER_134_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08974_ _15300_/Q _08981_/C _08913_/X vssd1 vssd1 vccd1 vccd1 _08976_/C sky130_fd_sc_hd__a21o_1
XFILLER_102_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_07925_ _09543_/A _07949_/B vssd1 vssd1 vccd1 vccd1 _07930_/A sky130_fd_sc_hd__xnor2_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07856_ _13824_/C _07989_/B vssd1 vssd1 vccd1 vccd1 _07857_/B sky130_fd_sc_hd__xnor2_4
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07787_ _15440_/Q _08144_/B vssd1 vssd1 vccd1 vccd1 _07828_/A sky130_fd_sc_hd__xnor2_4
X_09526_ _09524_/Y _09519_/C _09531_/A _09523_/Y vssd1 vssd1 vccd1 vccd1 _09531_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09457_ _09455_/Y _09449_/C _09451_/X _09454_/Y vssd1 vssd1 vccd1 vccd1 _09458_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08408_ _08414_/A _08414_/B vssd1 vssd1 vccd1 vccd1 _08468_/A sky130_fd_sc_hd__xor2_2
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09388_ _11229_/A vssd1 vssd1 vccd1 vccd1 _13532_/A sky130_fd_sc_hd__buf_4
XFILLER_8_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08339_ _08339_/A _08325_/A vssd1 vssd1 vccd1 vccd1 _08339_/X sky130_fd_sc_hd__or2b_1
X_11350_ _11343_/B _11344_/C _11347_/X _11348_/Y vssd1 vssd1 vccd1 vccd1 _11351_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10301_ _10301_/A _10301_/B _10301_/C vssd1 vssd1 vccd1 vccd1 _10302_/C sky130_fd_sc_hd__nand3_1
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11281_ _11373_/A _11281_/B _11286_/A vssd1 vssd1 vccd1 vccd1 _15657_/D sky130_fd_sc_hd__nor3_1
X_13020_ _13018_/Y _13014_/C _13025_/A _13017_/Y vssd1 vssd1 vccd1 vccd1 _13025_/B
+ sky130_fd_sc_hd__a211oi_1
X_10232_ _15502_/Q _15501_/Q _15500_/Q _10119_/X vssd1 vssd1 vccd1 vccd1 _15494_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10163_ _15484_/Q _10162_/C _10044_/X vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__a21oi_1
XFILLER_105_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10094_ _15472_/Q _10150_/B _10100_/C vssd1 vssd1 vccd1 vccd1 _10094_/Y sky130_fd_sc_hd__nand3_1
X_14971_ _14970_/X _14969_/A _14815_/X vssd1 vssd1 vccd1 vccd1 _14971_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13922_ _14316_/A vssd1 vssd1 vccd1 vccd1 _13922_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13853_ _16079_/Q _13853_/B _13853_/C vssd1 vssd1 vccd1 vccd1 _13861_/B sky130_fd_sc_hd__and3_1
XFILLER_90_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12804_ _12804_/A _12804_/B _12808_/B vssd1 vssd1 vccd1 vccd1 _15896_/D sky130_fd_sc_hd__nor3_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13784_ _13784_/A vssd1 vssd1 vccd1 vccd1 _16064_/D sky130_fd_sc_hd__clkbuf_1
X_10996_ _10996_/A _10996_/B _10996_/C vssd1 vssd1 vccd1 vccd1 _10997_/C sky130_fd_sc_hd__nand3_1
XFILLER_90_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15523_ _15655_/CLK _15523_/D vssd1 vssd1 vccd1 vccd1 _15523_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _15887_/Q _12954_/B _12742_/C vssd1 vssd1 vccd1 vccd1 _12735_/X sky130_fd_sc_hd__and3_1
XFILLER_43_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _15483_/CLK _15454_/D vssd1 vssd1 vccd1 vccd1 _15454_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12666_/A vssd1 vssd1 vccd1 vccd1 _15875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14405_ _14403_/X _14405_/B vssd1 vssd1 vccd1 vccd1 _14405_/X sky130_fd_sc_hd__and2b_1
X_11617_ _11653_/A _11617_/B _11617_/C vssd1 vssd1 vccd1 vccd1 _11618_/A sky130_fd_sc_hd__and3_1
X_15385_ _15484_/CLK _15385_/D vssd1 vssd1 vccd1 vccd1 _15385_/Q sky130_fd_sc_hd__dfxtp_1
X_12597_ _12598_/B _12598_/C _12598_/A vssd1 vssd1 vccd1 vccd1 _12599_/B sky130_fd_sc_hd__a21o_1
XFILLER_11_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14336_ _16174_/Q _14357_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14338_/B sky130_fd_sc_hd__a21oi_1
X_11548_ _15700_/Q _11547_/C _11488_/X vssd1 vssd1 vccd1 vccd1 _11549_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14267_ _14265_/A _14265_/B _14264_/Y _14266_/Y vssd1 vssd1 vccd1 vccd1 _16156_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_128_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ _15690_/Q _11655_/B _11479_/C vssd1 vssd1 vccd1 vccd1 _11491_/A sky130_fd_sc_hd__and3_1
X_13218_ _13218_/A _13218_/B _13222_/A vssd1 vssd1 vccd1 vccd1 _15964_/D sky130_fd_sc_hd__nor3_1
X_16006_ _16007_/CLK _16006_/D vssd1 vssd1 vccd1 vccd1 _16006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14198_ _14195_/X _14193_/B _14197_/Y vssd1 vssd1 vccd1 vccd1 _16141_/D sky130_fd_sc_hd__o21a_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13149_/A _13149_/B _13149_/C vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__and3_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _14970_/A vssd1 vssd1 vccd1 vccd1 _07710_/X sky130_fd_sc_hd__buf_2
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08690_ _08704_/A _08690_/B _08690_/C vssd1 vssd1 vccd1 vccd1 _08691_/A sky130_fd_sc_hd__and3_1
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07641_ input3/X vssd1 vssd1 vccd1 vccd1 _12661_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09311_ _15233_/Q _15232_/Q _15231_/Q _09194_/X vssd1 vssd1 vccd1 vccd1 _15351_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_34_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09242_ _15341_/Q _09354_/B _09242_/C vssd1 vssd1 vccd1 vccd1 _09251_/B sky130_fd_sc_hd__and3_1
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09173_ _15331_/Q _09290_/B _09173_/C vssd1 vssd1 vccd1 vccd1 _09183_/A sky130_fd_sc_hd__and3_1
X_08124_ _15223_/Q vssd1 vssd1 vccd1 vccd1 _09024_/A sky130_fd_sc_hd__clkinv_2
XFILLER_135_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08055_ _15719_/Q vssd1 vssd1 vccd1 vccd1 _11676_/A sky130_fd_sc_hd__inv_2
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ _08957_/A _08957_/B vssd1 vssd1 vccd1 vccd1 _08961_/C sky130_fd_sc_hd__nor2_1
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07908_ _07963_/B _07908_/B vssd1 vssd1 vccd1 vccd1 _07909_/B sky130_fd_sc_hd__nand2_4
X_08888_ _10044_/A vssd1 vssd1 vccd1 vccd1 _08888_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07839_ _15945_/Q vssd1 vssd1 vccd1 vccd1 _13162_/C sky130_fd_sc_hd__clkinv_2
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _15590_/Q _11023_/B _10855_/C vssd1 vssd1 vccd1 vccd1 _10850_/Y sky130_fd_sc_hd__nand3_1
XFILLER_112_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09509_ _09504_/X _09507_/Y _09508_/Y _09501_/C vssd1 vssd1 vccd1 vccd1 _09511_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ _10789_/A _10781_/B _10781_/C vssd1 vssd1 vccd1 vccd1 _10782_/A sky130_fd_sc_hd__and3_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12520_ _15853_/Q _12519_/C _12347_/X vssd1 vssd1 vccd1 vccd1 _12521_/B sky130_fd_sc_hd__a21oi_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _15841_/Q _12507_/B _12456_/C vssd1 vssd1 vccd1 vccd1 _12451_/Y sky130_fd_sc_hd__nand3_1
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11402_ _15678_/Q _11409_/C _11230_/X vssd1 vssd1 vccd1 vccd1 _11402_/Y sky130_fd_sc_hd__a21oi_1
X_15170_ _15170_/A vssd1 vssd1 vccd1 vccd1 _16361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12382_ _12382_/A vssd1 vssd1 vccd1 vccd1 _15830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14121_ _14122_/B _14122_/C _14122_/A vssd1 vssd1 vccd1 vccd1 _14123_/B sky130_fd_sc_hd__a21o_1
X_11333_ _11347_/C vssd1 vssd1 vccd1 vccd1 _11355_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14052_ _14045_/Y _14046_/X _14048_/B vssd1 vssd1 vccd1 vccd1 _14053_/B sky130_fd_sc_hd__o21a_1
X_11264_ _11264_/A _11264_/B vssd1 vssd1 vccd1 vccd1 _11268_/C sky130_fd_sc_hd__nor2_1
XFILLER_4_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13003_ _15931_/Q _13004_/C _13130_/A vssd1 vssd1 vccd1 vccd1 _13003_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10215_ _15492_/Q _10220_/C _09981_/X vssd1 vssd1 vccd1 vccd1 _10215_/Y sky130_fd_sc_hd__a21oi_1
X_11195_ _11193_/Y _11189_/C _11202_/A _11192_/Y vssd1 vssd1 vccd1 vccd1 _11202_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ _10153_/A _10146_/B _10146_/C vssd1 vssd1 vccd1 vccd1 _10147_/A sky130_fd_sc_hd__and3_1
XFILLER_79_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10077_ _10074_/X _10076_/Y _10071_/B _10072_/C vssd1 vssd1 vccd1 vccd1 _10079_/B
+ sky130_fd_sc_hd__o211ai_1
X_14954_ _16313_/Q _14953_/C _14917_/X vssd1 vssd1 vccd1 vccd1 _14955_/B sky130_fd_sc_hd__a21oi_1
X_13905_ _16088_/Q _13903_/C _15043_/A vssd1 vssd1 vccd1 vccd1 _13906_/B sky130_fd_sc_hd__a21o_1
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14885_ _15045_/A _14891_/C vssd1 vssd1 vccd1 vccd1 _14885_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13836_ _13844_/A _13836_/B _13836_/C vssd1 vssd1 vccd1 vccd1 _13837_/A sky130_fd_sc_hd__and3_1
XFILLER_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10979_ _11151_/A _10979_/B _10979_/C vssd1 vssd1 vccd1 vccd1 _10981_/B sky130_fd_sc_hd__or3_1
X_13767_ _13766_/B _13766_/C _13562_/X vssd1 vssd1 vccd1 vccd1 _13768_/C sky130_fd_sc_hd__o21ai_1
X_15506_ _15224_/Q _15506_/D vssd1 vssd1 vccd1 vccd1 _15506_/Q sky130_fd_sc_hd__dfxtp_1
X_12718_ _12740_/A _12718_/B _12718_/C vssd1 vssd1 vccd1 vccd1 _12719_/A sky130_fd_sc_hd__and3_1
X_13698_ _13735_/A _13698_/B _13698_/C vssd1 vssd1 vccd1 vccd1 _13699_/A sky130_fd_sc_hd__and3_1
X_15437_ _15484_/CLK _15437_/D vssd1 vssd1 vccd1 vccd1 _15437_/Q sky130_fd_sc_hd__dfxtp_1
X_12649_ _15874_/Q _12690_/C _12481_/X vssd1 vssd1 vccd1 vccd1 _12652_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15368_ _15368_/CLK _15368_/D vssd1 vssd1 vccd1 vccd1 _15368_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14319_ _14312_/Y _14313_/X _14315_/B vssd1 vssd1 vccd1 vccd1 _14320_/B sky130_fd_sc_hd__o21a_1
X_15299_ _16344_/CLK _15299_/D vssd1 vssd1 vccd1 vccd1 _15299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09860_ _15437_/Q _10029_/B _09867_/C vssd1 vssd1 vccd1 vccd1 _09860_/X sky130_fd_sc_hd__and3_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _15274_/Q _09047_/B _08811_/C vssd1 vssd1 vccd1 vccd1 _08811_/Y sky130_fd_sc_hd__nand3_1
X_09791_ _09791_/A vssd1 vssd1 vccd1 vccd1 _15425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08742_ _08742_/A _08742_/B _08742_/C vssd1 vssd1 vccd1 vccd1 _08743_/C sky130_fd_sc_hd__nand3_1
XFILLER_97_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08673_ _08686_/C vssd1 vssd1 vccd1 vccd1 _08694_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07624_ _15202_/Q _07658_/C _07623_/X vssd1 vssd1 vccd1 vccd1 _07626_/B sky130_fd_sc_hd__a21oi_1
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09225_ _09233_/A _09225_/B _09225_/C vssd1 vssd1 vccd1 vccd1 _09226_/A sky130_fd_sc_hd__and3_1
XFILLER_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09156_ _09171_/A _09156_/B _09156_/C vssd1 vssd1 vccd1 vccd1 _09157_/A sky130_fd_sc_hd__and3_1
X_08107_ _14941_/C _08107_/B vssd1 vssd1 vccd1 vccd1 _08107_/X sky130_fd_sc_hd__or2_1
XFILLER_108_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ _15317_/Q _09125_/C _09029_/X vssd1 vssd1 vccd1 vccd1 _09089_/B sky130_fd_sc_hd__a21oi_1
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08038_ _11275_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _08038_/X sky130_fd_sc_hd__or2_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10000_ _10000_/A vssd1 vssd1 vccd1 vccd1 _15457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09989_ _15457_/Q _10220_/B _09989_/C vssd1 vssd1 vccd1 vccd1 _09997_/B sky130_fd_sc_hd__and3_1
XFILLER_130_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11951_ _15763_/Q _11950_/C _11775_/X vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__a21oi_1
XFILLER_85_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10902_ _10902_/A _10902_/B _10902_/C vssd1 vssd1 vccd1 vccd1 _10903_/A sky130_fd_sc_hd__and3_1
XFILLER_45_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11882_ _11880_/Y _11875_/C _11878_/X _11879_/Y vssd1 vssd1 vccd1 vccd1 _11883_/C
+ sky130_fd_sc_hd__a211o_1
X_14670_ _14670_/A vssd1 vssd1 vccd1 vccd1 _16244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10833_ _10939_/C vssd1 vssd1 vccd1 vccd1 _12041_/A sky130_fd_sc_hd__buf_4
X_13621_ _13868_/A vssd1 vssd1 vccd1 vccd1 _13730_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater14 _15194_/Q vssd1 vssd1 vccd1 vccd1 _15655_/CLK sky130_fd_sc_hd__buf_12
X_16340_ _16359_/CLK _16340_/D vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
X_10764_ _15578_/Q _10876_/B _10770_/C vssd1 vssd1 vccd1 vccd1 _10767_/B sky130_fd_sc_hd__nand3_1
X_13552_ _13550_/Y _13546_/C _13557_/A _13549_/Y vssd1 vssd1 vccd1 vccd1 _13557_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12503_ _12510_/A _12503_/B _12503_/C vssd1 vssd1 vccd1 vccd1 _12504_/A sky130_fd_sc_hd__and3_1
X_16271_ _16273_/CLK _16271_/D vssd1 vssd1 vccd1 vccd1 _16271_/Q sky130_fd_sc_hd__dfxtp_2
X_13483_ _13612_/A vssd1 vssd1 vccd1 vccd1 _13538_/A sky130_fd_sc_hd__clkbuf_2
X_10695_ _10694_/B _10694_/C _10464_/X vssd1 vssd1 vccd1 vccd1 _10696_/C sky130_fd_sc_hd__o21ai_1
XFILLER_8_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15222_ _15254_/CLK _15222_/D vssd1 vssd1 vccd1 vccd1 state1[7] sky130_fd_sc_hd__dfxtp_2
X_12434_ _15840_/Q _12434_/B _12434_/C vssd1 vssd1 vccd1 vccd1 _12434_/X sky130_fd_sc_hd__and3_1
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15153_ _14408_/A _15155_/C _15086_/X vssd1 vssd1 vccd1 vccd1 _15154_/B sky130_fd_sc_hd__o21ai_1
X_12365_ _15829_/Q _12405_/C _12197_/X vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_101_clk _15665_/CLK vssd1 vssd1 vccd1 vccd1 _15728_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11316_ _11373_/A _11316_/B _11320_/B vssd1 vssd1 vccd1 vccd1 _15662_/D sky130_fd_sc_hd__nor3_1
X_14104_ _14644_/A _14106_/C vssd1 vssd1 vccd1 vccd1 _14104_/X sky130_fd_sc_hd__or2_1
X_15084_ _15084_/A _15084_/B vssd1 vssd1 vccd1 vccd1 _16338_/D sky130_fd_sc_hd__nor2_1
X_12296_ _12352_/A _12299_/C vssd1 vssd1 vccd1 vccd1 _12296_/X sky130_fd_sc_hd__or2_1
XFILLER_113_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14035_ _14040_/A _14034_/Y _14028_/B _14029_/C vssd1 vssd1 vccd1 vccd1 _14037_/B
+ sky130_fd_sc_hd__o211a_1
X_11247_ _11244_/X _11245_/Y _11246_/Y _11242_/C vssd1 vssd1 vccd1 vccd1 _11249_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_106_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11178_ _15642_/Q _11409_/B _11178_/C vssd1 vssd1 vccd1 vccd1 _11178_/Y sky130_fd_sc_hd__nand3_1
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10129_ _15479_/Q _10135_/C _10068_/X vssd1 vssd1 vccd1 vccd1 _10131_/C sky130_fd_sc_hd__a21o_1
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15986_ _16052_/CLK _15986_/D vssd1 vssd1 vccd1 vccd1 _15986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14937_ _14941_/C vssd1 vssd1 vccd1 vccd1 _14953_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14868_ _14868_/A vssd1 vssd1 vccd1 vccd1 _16289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13819_ _13824_/C vssd1 vssd1 vccd1 vccd1 _13832_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14799_ _14799_/A _14799_/B vssd1 vssd1 vccd1 vccd1 _14800_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09010_ _09018_/B _09010_/B vssd1 vssd1 vccd1 vccd1 _09012_/A sky130_fd_sc_hd__or2_1
XFILLER_148_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09912_ _09909_/X _09910_/Y _09911_/Y _09907_/C vssd1 vssd1 vccd1 vccd1 _09914_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _09843_/A _09843_/B _09843_/C vssd1 vssd1 vccd1 vccd1 _09844_/C sky130_fd_sc_hd__nand3_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _15424_/Q _09950_/B _09784_/C vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__and3_1
XFILLER_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08725_ _11037_/A vssd1 vssd1 vccd1 vccd1 _14372_/A sky130_fd_sc_hd__buf_4
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08656_ _08774_/A _08656_/B _08660_/B vssd1 vssd1 vccd1 vccd1 _15249_/D sky130_fd_sc_hd__nor3_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _13720_/A vssd1 vssd1 vccd1 vccd1 _09541_/A sky130_fd_sc_hd__buf_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08587_ _08611_/A _08587_/B _08593_/B vssd1 vssd1 vccd1 vccd1 _15240_/D sky130_fd_sc_hd__nor3_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09208_ _09208_/A _09208_/B _09208_/C vssd1 vssd1 vccd1 vccd1 _09209_/C sky130_fd_sc_hd__nand3_1
X_10480_ _10481_/B _10481_/C _10481_/A vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09139_ _09152_/C vssd1 vssd1 vccd1 vccd1 _09160_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12150_ _15795_/Q _12150_/B _12150_/C vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__and3_1
X_11101_ _11113_/C vssd1 vssd1 vccd1 vccd1 _11121_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12081_ _15784_/Q _12121_/C _11912_/X vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__a21oi_1
XFILLER_78_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ _11204_/A _11036_/C vssd1 vssd1 vccd1 vccd1 _11032_/X sky130_fd_sc_hd__or2_1
XFILLER_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15840_ _15907_/CLK _15840_/D vssd1 vssd1 vccd1 vccd1 _15840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15771_ _15195_/Q _15771_/D vssd1 vssd1 vccd1 vccd1 _15771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12983_ _12983_/A vssd1 vssd1 vccd1 vccd1 _12996_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14722_ _14722_/A _14722_/B vssd1 vssd1 vccd1 vccd1 _14723_/B sky130_fd_sc_hd__nor2_1
X_11934_ _11941_/A _11934_/B _11934_/C vssd1 vssd1 vccd1 vccd1 _11935_/A sky130_fd_sc_hd__and3_1
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14653_ _14653_/A vssd1 vssd1 vccd1 vccd1 _14811_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_11865_ _11863_/X _11864_/Y _11860_/B _11861_/C vssd1 vssd1 vccd1 vccd1 _11867_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_60_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13604_ _13604_/A _13604_/B _13608_/B vssd1 vssd1 vccd1 vccd1 _16031_/D sky130_fd_sc_hd__nor3_1
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10816_ _15586_/Q _10855_/C _10760_/X vssd1 vssd1 vccd1 vccd1 _10818_/B sky130_fd_sc_hd__a21oi_1
X_11796_ _11796_/A _11796_/B _11801_/A vssd1 vssd1 vccd1 vccd1 _15738_/D sky130_fd_sc_hd__nor3_1
X_14584_ _16228_/Q _15021_/A _14584_/C vssd1 vssd1 vccd1 vccd1 _14590_/A sky130_fd_sc_hd__and3_1
XFILLER_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16323_ _16359_/CLK _16323_/D vssd1 vssd1 vccd1 vccd1 _16323_/Q sky130_fd_sc_hd__dfxtp_1
X_13535_ _16022_/Q _13533_/C _13534_/X vssd1 vssd1 vccd1 vccd1 _13535_/Y sky130_fd_sc_hd__a21oi_1
X_10747_ _10745_/A _10745_/B _10746_/X vssd1 vssd1 vccd1 vccd1 _15573_/D sky130_fd_sc_hd__a21oi_1
XFILLER_146_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16254_ _16264_/CLK _16254_/D vssd1 vssd1 vccd1 vccd1 _16254_/Q sky130_fd_sc_hd__dfxtp_2
X_10678_ _11099_/A vssd1 vssd1 vccd1 vccd1 _10797_/A sky130_fd_sc_hd__buf_2
X_13466_ _13412_/X _13462_/C _13465_/Y vssd1 vssd1 vccd1 vccd1 _16007_/D sky130_fd_sc_hd__a21oi_1
X_15205_ _16241_/CLK _15205_/D vssd1 vssd1 vccd1 vccd1 _15205_/Q sky130_fd_sc_hd__dfxtp_1
X_12417_ _12417_/A vssd1 vssd1 vccd1 vccd1 _15835_/D sky130_fd_sc_hd__clkbuf_1
X_16185_ _16204_/CLK _16185_/D vssd1 vssd1 vccd1 vccd1 _16185_/Q sky130_fd_sc_hd__dfxtp_1
X_13397_ _13404_/A _13395_/Y _13396_/Y _13392_/C vssd1 vssd1 vccd1 vccd1 _13399_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15136_ _15136_/A vssd1 vssd1 vccd1 vccd1 _16352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ _15826_/Q _12346_/C _12347_/X vssd1 vssd1 vccd1 vccd1 _12349_/B sky130_fd_sc_hd__a21oi_1
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12279_ _12275_/X _12276_/Y _12278_/Y _12273_/C vssd1 vssd1 vccd1 vccd1 _12281_/B
+ sky130_fd_sc_hd__o211ai_1
X_15067_ _16339_/Q _15171_/B _15072_/C vssd1 vssd1 vccd1 vccd1 _15075_/A sky130_fd_sc_hd__and3_1
XFILLER_99_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14018_ _16232_/Q _16231_/Q _16230_/Q _13973_/X vssd1 vssd1 vccd1 vccd1 _16107_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15969_ _15970_/CLK _15969_/D vssd1 vssd1 vccd1 vccd1 _15969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08510_ input5/X vssd1 vssd1 vccd1 vccd1 _10896_/A sky130_fd_sc_hd__clkbuf_4
X_09490_ _09778_/A vssd1 vssd1 vccd1 vccd1 _09490_/X sky130_fd_sc_hd__buf_2
XFILLER_64_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08441_ _08442_/A _08442_/B vssd1 vssd1 vccd1 vccd1 _08443_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08372_ _08372_/A _08372_/B vssd1 vssd1 vccd1 vccd1 _08375_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09826_ _09997_/A _09826_/B _09826_/C vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__or3_1
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09757_ _09764_/B _09757_/B vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__or2_1
XFILLER_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _12616_/A vssd1 vssd1 vccd1 vccd1 _13700_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09685_/X _09686_/Y _09687_/Y _09683_/C vssd1 vssd1 vccd1 vccd1 _09690_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08648_/A _08639_/B _08639_/C vssd1 vssd1 vccd1 vccd1 _08640_/A sky130_fd_sc_hd__and3_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _15715_/Q _11650_/B _11655_/C vssd1 vssd1 vccd1 vccd1 _11650_/Y sky130_fd_sc_hd__nand3_1
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10601_ _10601_/A vssd1 vssd1 vccd1 vccd1 _15551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11581_ _11581_/A vssd1 vssd1 vccd1 vccd1 _15704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10532_ _15541_/Q _10532_/B _10540_/C vssd1 vssd1 vccd1 vccd1 _10537_/A sky130_fd_sc_hd__and3_1
X_13320_ _13348_/A _13320_/B _13324_/A vssd1 vssd1 vccd1 vccd1 _15982_/D sky130_fd_sc_hd__nor3_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10463_ _10577_/A _10463_/B _10463_/C vssd1 vssd1 vccd1 vccd1 _10466_/B sky130_fd_sc_hd__or3_1
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13251_ _14879_/A vssd1 vssd1 vccd1 vccd1 _13457_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12202_ _15803_/Q _12208_/C _12086_/X vssd1 vssd1 vccd1 vccd1 _12204_/C sky130_fd_sc_hd__a21o_1
XFILLER_129_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13182_ _13178_/X _13180_/Y _13181_/Y _13176_/C vssd1 vssd1 vccd1 vccd1 _13184_/B
+ sky130_fd_sc_hd__o211ai_1
X_10394_ _10511_/A _10394_/B _10398_/B vssd1 vssd1 vccd1 vccd1 _15518_/D sky130_fd_sc_hd__nor3_1
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12133_ _12133_/A vssd1 vssd1 vccd1 vccd1 _15790_/D sky130_fd_sc_hd__clkbuf_1
X_12064_ _15781_/Q _12062_/C _12063_/X vssd1 vssd1 vccd1 vccd1 _12065_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11015_ _15617_/Q _11021_/C _10897_/X vssd1 vssd1 vccd1 vccd1 _11015_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_104_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15823_ _15907_/CLK _15823_/D vssd1 vssd1 vccd1 vccd1 _15823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15754_ _15763_/CLK _15754_/D vssd1 vssd1 vccd1 vccd1 _15754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12966_ _12964_/Y _12959_/C _12971_/A _12963_/Y vssd1 vssd1 vccd1 vccd1 _12971_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14705_ _14716_/A _14705_/B _14709_/A vssd1 vssd1 vccd1 vccd1 _16252_/D sky130_fd_sc_hd__nor3_1
X_11917_ _15758_/Q _11923_/C _11798_/X vssd1 vssd1 vccd1 vccd1 _11919_/C sky130_fd_sc_hd__a21o_1
X_15685_ _15763_/CLK _15685_/D vssd1 vssd1 vccd1 vccd1 _15685_/Q sky130_fd_sc_hd__dfxtp_1
X_12897_ _12893_/X _12894_/Y _12896_/Y _12891_/C vssd1 vssd1 vccd1 vccd1 _12899_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_61_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14636_ _14642_/A _14635_/Y _14630_/B _14631_/C vssd1 vssd1 vccd1 vccd1 _14638_/B
+ sky130_fd_sc_hd__o211a_1
X_11848_ _15754_/Q _15753_/Q _15752_/Q _11847_/X vssd1 vssd1 vccd1 vccd1 _15746_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14567_ _16223_/Q _14566_/C _07674_/A vssd1 vssd1 vccd1 vccd1 _14568_/B sky130_fd_sc_hd__a21o_1
X_11779_ _11779_/A _11779_/B vssd1 vssd1 vccd1 vccd1 _11784_/C sky130_fd_sc_hd__nor2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16306_ _16317_/CLK _16306_/D vssd1 vssd1 vccd1 vccd1 _16306_/Q sky130_fd_sc_hd__dfxtp_2
X_13518_ _16034_/Q _16033_/Q _16032_/Q _13467_/X vssd1 vssd1 vccd1 vccd1 _16017_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_146_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14498_ _14328_/X _14372_/X _14493_/B _14459_/X vssd1 vssd1 vccd1 vccd1 _14499_/B
+ sky130_fd_sc_hd__a31o_1
X_16237_ _16247_/CLK _16237_/D vssd1 vssd1 vccd1 vccd1 _16237_/Q sky130_fd_sc_hd__dfxtp_2
X_13449_ _13447_/Y _13442_/C _13455_/A _13446_/Y vssd1 vssd1 vccd1 vccd1 _13455_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16168_ _16169_/CLK _16168_/D vssd1 vssd1 vccd1 vccd1 _16168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15119_ _15119_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _16347_/D sky130_fd_sc_hd__nor2_1
XFILLER_141_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08990_ _08987_/X _08988_/Y _08989_/Y _08985_/C vssd1 vssd1 vccd1 vccd1 _08992_/B
+ sky130_fd_sc_hd__o211ai_1
X_16099_ _16100_/CLK _16099_/D vssd1 vssd1 vccd1 vccd1 _16099_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07941_ _08610_/C vssd1 vssd1 vccd1 vccd1 _08622_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07872_ _16071_/Q _16089_/Q vssd1 vssd1 vccd1 vccd1 _07873_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09611_ _09612_/B _09612_/C _09612_/A vssd1 vssd1 vccd1 vccd1 _09613_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09542_ _15394_/Q _15393_/Q _15392_/Q _09541_/X vssd1 vssd1 vccd1 vccd1 _15386_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09473_ _09471_/A _09471_/B _09472_/X vssd1 vssd1 vccd1 vccd1 _15375_/D sky130_fd_sc_hd__a21oi_1
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08424_ _08429_/C _08424_/B vssd1 vssd1 vccd1 vccd1 _08424_/Y sky130_fd_sc_hd__xnor2_1
X_08355_ _08356_/A _08356_/B _08356_/C vssd1 vssd1 vccd1 vccd1 _08388_/A sky130_fd_sc_hd__a21oi_4
XFILLER_149_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08286_ _08199_/A _08199_/B _08285_/X vssd1 vssd1 vccd1 vccd1 _08325_/A sky130_fd_sc_hd__a21bo_2
XFILLER_50_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09809_ _11963_/A vssd1 vssd1 vccd1 vccd1 _10388_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12820_ _12832_/C vssd1 vssd1 vccd1 vccd1 _12840_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12751_/A _12751_/B vssd1 vssd1 vccd1 vccd1 _12752_/B sky130_fd_sc_hd__nor2_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15422_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _15725_/Q _11819_/B _11712_/C vssd1 vssd1 vccd1 vccd1 _11702_/X sky130_fd_sc_hd__and3_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15470_ _15483_/CLK _15470_/D vssd1 vssd1 vccd1 vccd1 _15470_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _14541_/A vssd1 vssd1 vccd1 vccd1 _13239_/A sky130_fd_sc_hd__buf_2
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14421_ _14818_/A vssd1 vssd1 vccd1 vccd1 _14421_/X sky130_fd_sc_hd__clkbuf_4
X_11633_ _11633_/A vssd1 vssd1 vccd1 vccd1 _15712_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14352_ _14352_/A _14352_/B vssd1 vssd1 vccd1 vccd1 _14352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11564_ _11585_/C vssd1 vssd1 vccd1 vccd1 _11599_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _13301_/A _13301_/B _13302_/X vssd1 vssd1 vccd1 vccd1 _15978_/D sky130_fd_sc_hd__a21oi_1
X_10515_ _10515_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10516_/B sky130_fd_sc_hd__nor2_1
X_11495_ _11555_/A vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14283_ _14283_/A _14283_/B vssd1 vssd1 vccd1 vccd1 _16160_/D sky130_fd_sc_hd__nor2_1
XFILLER_109_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16022_ _16022_/CLK _16022_/D vssd1 vssd1 vccd1 vccd1 _16022_/Q sky130_fd_sc_hd__dfxtp_1
X_10446_ _15528_/Q _10446_/B _10446_/C vssd1 vssd1 vccd1 vccd1 _10456_/A sky130_fd_sc_hd__and3_1
X_13234_ _15968_/Q _13286_/B _13240_/C vssd1 vssd1 vccd1 vccd1 _13234_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10377_ _10375_/Y _10368_/C _10372_/X _10374_/Y vssd1 vssd1 vccd1 vccd1 _10378_/C
+ sky130_fd_sc_hd__a211o_1
X_13165_ _13679_/A vssd1 vssd1 vccd1 vccd1 _13374_/B sky130_fd_sc_hd__buf_2
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12116_ _15789_/Q _12121_/C _12001_/X vssd1 vssd1 vccd1 vccd1 _12116_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13096_ _13474_/A vssd1 vssd1 vccd1 vccd1 _14379_/A sky130_fd_sc_hd__clkbuf_4
X_12047_ _15779_/Q _12107_/B _12055_/C vssd1 vssd1 vccd1 vccd1 _12047_/X sky130_fd_sc_hd__and3_1
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15806_ _07603_/A _15806_/D vssd1 vssd1 vccd1 vccd1 _15806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13998_ _13998_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15737_ _15746_/CLK _15737_/D vssd1 vssd1 vccd1 vccd1 _15737_/Q sky130_fd_sc_hd__dfxtp_2
X_12949_ _15921_/Q _14031_/A _12949_/C vssd1 vssd1 vccd1 vccd1 _12949_/Y sky130_fd_sc_hd__nand3_1
XFILLER_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15312_/CLK sky130_fd_sc_hd__clkbuf_16
X_15668_ _15763_/CLK _15668_/D vssd1 vssd1 vccd1 vccd1 _15668_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_14619_ _14619_/A _14619_/B vssd1 vssd1 vccd1 vccd1 _16232_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15599_ _15194_/Q _15599_/D vssd1 vssd1 vccd1 vccd1 _15599_/Q sky130_fd_sc_hd__dfxtp_1
X_08140_ _15548_/Q _08140_/B vssd1 vssd1 vccd1 vccd1 _08140_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08071_ _15665_/Q vssd1 vssd1 vccd1 vccd1 _11332_/A sky130_fd_sc_hd__inv_2
XFILLER_119_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08973_ _15300_/Q _09146_/B _08981_/C vssd1 vssd1 vccd1 vccd1 _08976_/B sky130_fd_sc_hd__nand3_1
XFILLER_102_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07924_ _10002_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07949_/B sky130_fd_sc_hd__xnor2_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07855_ _16161_/Q _07996_/B vssd1 vssd1 vccd1 vccd1 _07989_/B sky130_fd_sc_hd__xnor2_2
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07786_ _07786_/A _07786_/B vssd1 vssd1 vccd1 vccd1 _08144_/B sky130_fd_sc_hd__xor2_4
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09525_ _09531_/A _09523_/Y _09524_/Y _09519_/C vssd1 vssd1 vccd1 vccd1 _09527_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _16352_/CLK sky130_fd_sc_hd__clkbuf_16
X_09456_ _09451_/X _09454_/Y _09455_/Y _09449_/C vssd1 vssd1 vccd1 vccd1 _09458_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _08388_/A _08388_/B _08406_/X vssd1 vssd1 vccd1 vccd1 _08414_/B sky130_fd_sc_hd__a21oi_2
X_09387_ _15364_/Q _09391_/C _09220_/X vssd1 vssd1 vccd1 vccd1 _09387_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08338_ _08326_/B _08338_/B vssd1 vssd1 vccd1 vccd1 _08391_/A sky130_fd_sc_hd__and2b_2
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08269_ _08270_/A _08270_/B _08270_/C vssd1 vssd1 vccd1 vccd1 _08271_/A sky130_fd_sc_hd__a21oi_2
XFILLER_125_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10300_ _10301_/B _10301_/C _10301_/A vssd1 vssd1 vccd1 vccd1 _10302_/B sky130_fd_sc_hd__a21o_1
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11280_ _15658_/Q _11449_/B _11289_/C vssd1 vssd1 vccd1 vccd1 _11286_/A sky130_fd_sc_hd__and3_1
XFILLER_137_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10231_ _10231_/A vssd1 vssd1 vccd1 vccd1 _15493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10162_ _15484_/Q _10220_/B _10162_/C vssd1 vssd1 vccd1 vccd1 _10171_/B sky130_fd_sc_hd__and3_1
XFILLER_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10093_ _15473_/Q _10100_/C _10030_/X vssd1 vssd1 vccd1 vccd1 _10093_/Y sky130_fd_sc_hd__a21oi_1
X_14970_ _14970_/A vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13921_ _14325_/A vssd1 vssd1 vccd1 vccd1 _13921_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13852_ _13852_/A _13852_/B _13856_/B vssd1 vssd1 vccd1 vccd1 _16076_/D sky130_fd_sc_hd__nor3_1
X_12803_ _12801_/Y _12796_/C _12808_/A _12799_/Y vssd1 vssd1 vccd1 vccd1 _12808_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13783_ _13789_/A _13783_/B _13783_/C vssd1 vssd1 vccd1 vccd1 _13784_/A sky130_fd_sc_hd__and3_1
X_10995_ _10996_/B _10996_/C _10996_/A vssd1 vssd1 vccd1 vccd1 _10997_/B sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_54_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16304_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15522_ _15655_/CLK _15522_/D vssd1 vssd1 vccd1 vccd1 _15522_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12734_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12954_/B sky130_fd_sc_hd__buf_2
XFILLER_35_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15453_ _15483_/CLK _15453_/D vssd1 vssd1 vccd1 vccd1 _15453_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12680_/A _12665_/B _12665_/C vssd1 vssd1 vccd1 vccd1 _12666_/A sky130_fd_sc_hd__and3_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _16187_/Q _14403_/C _14270_/X vssd1 vssd1 vccd1 vccd1 _14405_/B sky130_fd_sc_hd__a21o_1
X_11616_ _11614_/B _11614_/C _11615_/X vssd1 vssd1 vccd1 vccd1 _11617_/C sky130_fd_sc_hd__o21ai_1
X_15384_ _15484_/CLK _15384_/D vssd1 vssd1 vccd1 vccd1 _15384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12596_ _15866_/Q _12601_/C _12370_/X vssd1 vssd1 vccd1 vccd1 _12598_/C sky130_fd_sc_hd__a21o_1
XFILLER_128_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14335_ _14345_/C vssd1 vssd1 vccd1 vccd1 _14357_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11547_ _15700_/Q _11719_/B _11547_/C vssd1 vssd1 vccd1 vccd1 _11556_/B sky130_fd_sc_hd__and3_1
XFILLER_144_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14266_ _14265_/X _14264_/Y _14042_/X vssd1 vssd1 vccd1 vccd1 _14266_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11478_ _11478_/A vssd1 vssd1 vccd1 vccd1 _15688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16005_ _16007_/CLK _16005_/D vssd1 vssd1 vccd1 vccd1 _16005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13217_ _15966_/Q _13420_/B _13217_/C vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__and3_1
X_10429_ _10421_/B _10422_/C _10426_/X _10427_/Y vssd1 vssd1 vccd1 vccd1 _10430_/C
+ sky130_fd_sc_hd__a211o_1
X_14197_ _14149_/X _14193_/B _14196_/X vssd1 vssd1 vccd1 vccd1 _14197_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13148_ _13146_/B _13146_/C _14892_/A vssd1 vssd1 vccd1 vccd1 _13149_/C sky130_fd_sc_hd__o21ai_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _15944_/Q _13078_/C _10970_/C vssd1 vssd1 vccd1 vccd1 _13080_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ _07640_/A vssd1 vssd1 vccd1 vccd1 _15199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_45_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16240_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09310_ _09310_/A vssd1 vssd1 vccd1 vccd1 _15350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ _09353_/A _09241_/B _09245_/B vssd1 vssd1 vccd1 vccd1 _15339_/D sky130_fd_sc_hd__nor3_1
X_09172_ _09172_/A vssd1 vssd1 vccd1 vccd1 _15329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08123_ _15225_/Q vssd1 vssd1 vccd1 vccd1 _08546_/A sky130_fd_sc_hd__inv_2
XFILLER_147_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _15701_/Q vssd1 vssd1 vccd1 vccd1 _11562_/A sky130_fd_sc_hd__inv_2
XFILLER_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08956_ _10110_/A vssd1 vssd1 vccd1 vccd1 _09185_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07907_ _07963_/A _07906_/C _16269_/Q vssd1 vssd1 vccd1 vccd1 _07908_/B sky130_fd_sc_hd__a21o_1
X_08887_ _10969_/A vssd1 vssd1 vccd1 vccd1 _10044_/A sky130_fd_sc_hd__buf_4
XFILLER_57_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07838_ _14207_/C _08025_/B vssd1 vssd1 vccd1 vccd1 _07844_/A sky130_fd_sc_hd__xnor2_4
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07769_ _15611_/Q _15593_/Q vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_36_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16362_/CLK sky130_fd_sc_hd__clkbuf_16
X_09508_ _15381_/Q _09623_/B _09508_/C vssd1 vssd1 vccd1 vccd1 _09508_/Y sky130_fd_sc_hd__nand3_1
XFILLER_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10778_/Y _10774_/C _10776_/X _10777_/Y vssd1 vssd1 vccd1 vccd1 _10781_/C
+ sky130_fd_sc_hd__a211o_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _15372_/Q _09446_/C _09212_/X vssd1 vssd1 vccd1 vccd1 _09439_/Y sky130_fd_sc_hd__a21oi_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _15842_/Q _12456_/C _12332_/X vssd1 vssd1 vccd1 vccd1 _12450_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _15678_/Q _11576_/B _11401_/C vssd1 vssd1 vccd1 vccd1 _11401_/X sky130_fd_sc_hd__and3_1
X_12381_ _12396_/A _12381_/B _12381_/C vssd1 vssd1 vccd1 vccd1 _12382_/A sky130_fd_sc_hd__and3_1
XFILLER_126_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14120_ _16130_/Q _14125_/C _13982_/X vssd1 vssd1 vccd1 vccd1 _14122_/C sky130_fd_sc_hd__a21o_1
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ _11332_/A vssd1 vssd1 vccd1 vccd1 _11347_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14051_ _14045_/Y _14048_/X _14050_/Y vssd1 vssd1 vccd1 vccd1 _16112_/D sky130_fd_sc_hd__o21a_1
XFILLER_125_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11263_ _11551_/A vssd1 vssd1 vccd1 vccd1 _11493_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13002_ _15931_/Q _13057_/B _13004_/C vssd1 vssd1 vccd1 vccd1 _13002_/X sky130_fd_sc_hd__and3_1
X_10214_ _15492_/Q _10446_/B _10214_/C vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__and3_1
X_11194_ _11202_/A _11192_/Y _11193_/Y _11189_/C vssd1 vssd1 vccd1 vccd1 _11196_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10145_ _10143_/Y _10139_/C _10141_/X _10142_/Y vssd1 vssd1 vccd1 vccd1 _10146_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_94_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10076_ _15471_/Q _10085_/C _10075_/X vssd1 vssd1 vccd1 vccd1 _10076_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14953_ _16313_/Q _14953_/B _14953_/C vssd1 vssd1 vccd1 vccd1 _14955_/A sky130_fd_sc_hd__and3_1
X_13904_ _14270_/A vssd1 vssd1 vccd1 vccd1 _15043_/A sky130_fd_sc_hd__buf_2
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14884_ _14877_/A _14881_/B _14845_/X vssd1 vssd1 vccd1 vccd1 _14891_/C sky130_fd_sc_hd__o21a_1
XFILLER_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13835_ _13829_/B _13830_/C _13832_/X _13833_/Y vssd1 vssd1 vccd1 vccd1 _13836_/C
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_27_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _16123_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13766_ _14106_/A _13766_/B _13766_/C vssd1 vssd1 vccd1 vccd1 _13768_/B sky130_fd_sc_hd__or3_1
X_10978_ _10978_/A vssd1 vssd1 vccd1 vccd1 _11019_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _15224_/Q _15505_/D vssd1 vssd1 vccd1 vccd1 _15505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ _12717_/A _12717_/B _12717_/C vssd1 vssd1 vccd1 vccd1 _12718_/C sky130_fd_sc_hd__nand3_1
X_13697_ _13695_/Y _13690_/C _13692_/X _13694_/Y vssd1 vssd1 vccd1 vccd1 _13698_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15436_ _15483_/CLK _15436_/D vssd1 vssd1 vccd1 vccd1 _15436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _12684_/C vssd1 vssd1 vccd1 vccd1 _12690_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15367_ _15440_/CLK _15367_/D vssd1 vssd1 vccd1 vccd1 _15367_/Q sky130_fd_sc_hd__dfxtp_1
X_12579_ _12579_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _12583_/C sky130_fd_sc_hd__nor2_1
XFILLER_144_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14318_ _14312_/Y _14315_/X _14317_/Y vssd1 vssd1 vccd1 vccd1 _16166_/D sky130_fd_sc_hd__o21a_1
XFILLER_116_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15298_ _16344_/CLK _15298_/D vssd1 vssd1 vccd1 vccd1 _15298_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14249_ _16157_/Q _14249_/B _14256_/C vssd1 vssd1 vccd1 vccd1 _14253_/B sky130_fd_sc_hd__nand3_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _13534_/A vssd1 vssd1 vccd1 vccd1 _09047_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_112_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09807_/A _09790_/B _09790_/C vssd1 vssd1 vccd1 vccd1 _09791_/A sky130_fd_sc_hd__and3_1
XFILLER_85_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _08742_/B _08742_/C _08742_/A vssd1 vssd1 vccd1 vccd1 _08743_/B sky130_fd_sc_hd__a21o_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08672_ _15243_/Q vssd1 vssd1 vccd1 vccd1 _08686_/C sky130_fd_sc_hd__inv_2
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07623_ _08735_/A vssd1 vssd1 vccd1 vccd1 _07623_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _16052_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _09222_/Y _09216_/C _09219_/X _09221_/Y vssd1 vssd1 vccd1 vccd1 _09225_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09155_ _09149_/B _09150_/C _09152_/X _09153_/Y vssd1 vssd1 vccd1 vccd1 _09156_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08106_ _08106_/A vssd1 vssd1 vccd1 vccd1 _14941_/C sky130_fd_sc_hd__buf_2
X_09086_ _09117_/C vssd1 vssd1 vccd1 vccd1 _09125_/C sky130_fd_sc_hd__clkbuf_2
X_08037_ _08037_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__xnor2_4
XFILLER_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09988_ _11197_/A vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08939_ _15293_/Q _08996_/B _08945_/C vssd1 vssd1 vccd1 vccd1 _08939_/Y sky130_fd_sc_hd__nand3_1
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11950_ _15763_/Q _12007_/B _11950_/C vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__and3_1
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10901_ _10899_/Y _10893_/C _10895_/X _10898_/Y vssd1 vssd1 vccd1 vccd1 _10902_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_57_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11881_ _11878_/X _11879_/Y _11880_/Y _11875_/C vssd1 vssd1 vccd1 vccd1 _11883_/B
+ sky130_fd_sc_hd__o211ai_1
X_13620_ _16052_/Q _16051_/Q _16050_/Q _13467_/X vssd1 vssd1 vccd1 vccd1 _16035_/D
+ sky130_fd_sc_hd__o31a_1
X_10832_ _15589_/Q _10835_/C _10663_/X vssd1 vssd1 vccd1 vccd1 _10832_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater15 _15484_/CLK vssd1 vssd1 vccd1 vccd1 _15483_/CLK sky130_fd_sc_hd__buf_12
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13551_ _13557_/A _13549_/Y _13550_/Y _13546_/C vssd1 vssd1 vccd1 vccd1 _13553_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10763_ _10797_/A _10763_/B _10767_/A vssd1 vssd1 vccd1 vccd1 _15576_/D sky130_fd_sc_hd__nor3_1
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ _12500_/Y _12496_/C _12498_/X _12499_/Y vssd1 vssd1 vccd1 vccd1 _12503_/C
+ sky130_fd_sc_hd__a211o_1
X_16270_ _16273_/CLK _16270_/D vssd1 vssd1 vccd1 vccd1 _16270_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13482_ _13482_/A vssd1 vssd1 vccd1 vccd1 _16010_/D sky130_fd_sc_hd__clkbuf_1
X_10694_ _10863_/A _10694_/B _10694_/C vssd1 vssd1 vccd1 vccd1 _10696_/B sky130_fd_sc_hd__or3_1
XFILLER_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15221_ _16242_/CLK _15221_/D vssd1 vssd1 vccd1 vccd1 state1[6] sky130_fd_sc_hd__dfxtp_4
X_12433_ _12433_/A vssd1 vssd1 vccd1 vccd1 _15838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15152_ _15152_/A _15155_/C vssd1 vssd1 vccd1 vccd1 _15154_/A sky130_fd_sc_hd__and2_1
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12364_ _12399_/C vssd1 vssd1 vccd1 vccd1 _12405_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14103_ _14103_/A _14103_/B vssd1 vssd1 vccd1 vccd1 _14106_/C sky130_fd_sc_hd__nor2_1
X_11315_ _11313_/Y _11309_/C _11320_/A _11312_/Y vssd1 vssd1 vccd1 vccd1 _11320_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15083_ _14964_/X _15085_/C _15007_/X vssd1 vssd1 vccd1 vccd1 _15084_/B sky130_fd_sc_hd__o21ai_1
X_12295_ _12295_/A _12295_/B vssd1 vssd1 vccd1 vccd1 _12299_/C sky130_fd_sc_hd__nor2_1
XFILLER_107_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14034_ _16113_/Q _14032_/C _14033_/X vssd1 vssd1 vccd1 vccd1 _14034_/Y sky130_fd_sc_hd__a21oi_1
X_11246_ _15652_/Q _11362_/B _11253_/C vssd1 vssd1 vccd1 vccd1 _11246_/Y sky130_fd_sc_hd__nand3_1
XFILLER_122_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11177_ _12041_/A vssd1 vssd1 vccd1 vccd1 _11409_/B sky130_fd_sc_hd__buf_2
X_10128_ _15479_/Q _10298_/B _10135_/C vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__nand3_1
XFILLER_95_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15985_ _15994_/CLK _15985_/D vssd1 vssd1 vccd1 vccd1 _15985_/Q sky130_fd_sc_hd__dfxtp_1
X_10059_ _10074_/C vssd1 vssd1 vccd1 vccd1 _10085_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14936_ _14936_/A vssd1 vssd1 vccd1 vccd1 _15023_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14867_ _14946_/A _14867_/B _14867_/C vssd1 vssd1 vccd1 vccd1 _14868_/A sky130_fd_sc_hd__and3_1
XFILLER_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13818_ _16124_/Q _16123_/Q _16122_/Q _13723_/X vssd1 vssd1 vccd1 vccd1 _16071_/D
+ sky130_fd_sc_hd__o31a_1
X_14798_ _14798_/A _14798_/B vssd1 vssd1 vccd1 vccd1 _14799_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13749_ _13789_/A _13749_/B _13749_/C vssd1 vssd1 vccd1 vccd1 _13750_/A sky130_fd_sc_hd__and3_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15419_ _15484_/CLK _15419_/D vssd1 vssd1 vccd1 vccd1 _15419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15899_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09911_ _15444_/Q _09911_/B _09911_/C vssd1 vssd1 vccd1 vccd1 _09911_/Y sky130_fd_sc_hd__nand3_1
XFILLER_104_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _09843_/B _09843_/C _09843_/A vssd1 vssd1 vccd1 vccd1 _09844_/B sky130_fd_sc_hd__a21o_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _15424_/Q _09817_/C _09605_/X vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__a21oi_1
XFILLER_100_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08724_ _08839_/A _08724_/B _08724_/C vssd1 vssd1 vccd1 vccd1 _08728_/B sky130_fd_sc_hd__or3_1
XFILLER_73_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _08653_/Y _08648_/C _08660_/A _08652_/Y vssd1 vssd1 vccd1 vccd1 _08660_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _08722_/A vssd1 vssd1 vccd1 vccd1 _13720_/A sky130_fd_sc_hd__buf_8
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08586_ _08584_/Y _08580_/C _08593_/A _08583_/Y vssd1 vssd1 vccd1 vccd1 _08593_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_54_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09207_ _09208_/B _09208_/C _09208_/A vssd1 vssd1 vccd1 vccd1 _09209_/B sky130_fd_sc_hd__a21o_1
XFILLER_139_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09138_ _09138_/A vssd1 vssd1 vccd1 vccd1 _09152_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09069_ _09075_/B _09069_/B vssd1 vssd1 vccd1 vccd1 _09071_/A sky130_fd_sc_hd__or2_1
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11100_ _15629_/Q vssd1 vssd1 vccd1 vccd1 _11113_/C sky130_fd_sc_hd__inv_2
XFILLER_135_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12080_ _12115_/C vssd1 vssd1 vccd1 vccd1 _12121_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _11031_/A _11031_/B vssd1 vssd1 vccd1 vccd1 _11036_/C sky130_fd_sc_hd__nor2_1
XFILLER_89_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15770_ _15794_/CLK _15770_/D vssd1 vssd1 vccd1 vccd1 _15770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12982_ _15932_/Q _15934_/Q _15933_/Q _12981_/X vssd1 vssd1 vccd1 vccd1 _15926_/D
+ sky130_fd_sc_hd__o31a_1
X_14721_ _14721_/A _14721_/B vssd1 vssd1 vccd1 vccd1 _14722_/B sky130_fd_sc_hd__nor2_1
X_11933_ _11931_/Y _11927_/C _11929_/X _11930_/Y vssd1 vssd1 vccd1 vccd1 _11934_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ _14652_/A _14652_/B vssd1 vssd1 vccd1 vccd1 _16239_/D sky130_fd_sc_hd__nor2_1
X_11864_ _15750_/Q _11872_/C _11805_/X vssd1 vssd1 vccd1 vccd1 _11864_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13603_ _13601_/Y _13595_/C _13608_/A _13599_/Y vssd1 vssd1 vccd1 vccd1 _13608_/B
+ sky130_fd_sc_hd__a211oi_1
X_10815_ _10847_/C vssd1 vssd1 vccd1 vccd1 _10855_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14583_ _16228_/Q _14605_/C _14503_/X vssd1 vssd1 vccd1 vccd1 _14585_/B sky130_fd_sc_hd__a21oi_1
X_11795_ _15739_/Q _12025_/B _11804_/C vssd1 vssd1 vccd1 vccd1 _11801_/A sky130_fd_sc_hd__and3_1
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16322_ _16359_/CLK _16322_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
X_13534_ _13534_/A vssd1 vssd1 vccd1 vccd1 _13534_/X sky130_fd_sc_hd__clkbuf_4
X_10746_ _10916_/A _10750_/C vssd1 vssd1 vccd1 vccd1 _10746_/X sky130_fd_sc_hd__or2_1
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16253_ _16264_/CLK _16253_/D vssd1 vssd1 vccd1 vccd1 _16253_/Q sky130_fd_sc_hd__dfxtp_2
X_13465_ _13362_/X _13462_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13465_/Y sky130_fd_sc_hd__o21ai_1
X_10677_ _10677_/A vssd1 vssd1 vccd1 vccd1 _15562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ _16241_/CLK _15204_/D vssd1 vssd1 vccd1 vccd1 _15204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12416_ _12454_/A _12416_/B _12416_/C vssd1 vssd1 vccd1 vccd1 _12417_/A sky130_fd_sc_hd__and3_1
X_16184_ _16192_/CLK _16184_/D vssd1 vssd1 vccd1 vccd1 _16184_/Q sky130_fd_sc_hd__dfxtp_1
X_13396_ _15996_/Q _13550_/B _13401_/C vssd1 vssd1 vccd1 vccd1 _13396_/Y sky130_fd_sc_hd__nand3_1
X_15135_ _15135_/A _15135_/B _15135_/C vssd1 vssd1 vccd1 vccd1 _15136_/A sky130_fd_sc_hd__and3_1
XFILLER_127_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12347_ _12631_/A vssd1 vssd1 vccd1 vccd1 _12347_/X sky130_fd_sc_hd__buf_2
XFILLER_142_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15066_ _15066_/A vssd1 vssd1 vccd1 vccd1 _16334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12278_ _15814_/Q _12507_/B _12284_/C vssd1 vssd1 vccd1 vccd1 _12278_/Y sky130_fd_sc_hd__nand3_1
XFILLER_141_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14017_ _14017_/A _14017_/B vssd1 vssd1 vccd1 vccd1 _16106_/D sky130_fd_sc_hd__nor2_1
XFILLER_141_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11229_ _11229_/A vssd1 vssd1 vccd1 vccd1 _12377_/A sky130_fd_sc_hd__buf_4
XFILLER_110_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15968_ _15970_/CLK _15968_/D vssd1 vssd1 vccd1 vccd1 _15968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14919_ _14919_/A _14919_/B vssd1 vssd1 vccd1 vccd1 _14921_/A sky130_fd_sc_hd__or2_1
X_15899_ _15899_/CLK _15899_/D vssd1 vssd1 vccd1 vccd1 _15899_/Q sky130_fd_sc_hd__dfxtp_2
X_08440_ state1[5] _08462_/B vssd1 vssd1 vccd1 vccd1 _08442_/B sky130_fd_sc_hd__and2_1
XFILLER_17_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08371_ _08442_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08372_/B sky130_fd_sc_hd__or2_1
XFILLER_118_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09825_ _09825_/A vssd1 vssd1 vccd1 vccd1 _09865_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09756_ _15421_/Q _09754_/C _09755_/X vssd1 vssd1 vccd1 vccd1 _09757_/B sky130_fd_sc_hd__a21oi_1
XFILLER_101_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08707_ _15259_/Q _08715_/C _08524_/X vssd1 vssd1 vccd1 vccd1 _08707_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _15409_/Q _09862_/B _09692_/C vssd1 vssd1 vccd1 vccd1 _09687_/Y sky130_fd_sc_hd__nand3_1
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _08636_/Y _08629_/C _08632_/X _08635_/Y vssd1 vssd1 vccd1 vccd1 _08639_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _08566_/X _08567_/Y _08568_/Y _08564_/C vssd1 vssd1 vccd1 vccd1 _08571_/B
+ sky130_fd_sc_hd__o211ai_1
X_10600_ _10615_/A _10600_/B _10600_/C vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__and3_1
XFILLER_23_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11580_ _11597_/A _11580_/B _11580_/C vssd1 vssd1 vccd1 vccd1 _11581_/A sky130_fd_sc_hd__and3_1
XFILLER_128_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10531_ _15541_/Q _10569_/C _10474_/X vssd1 vssd1 vccd1 vccd1 _10533_/B sky130_fd_sc_hd__a21oi_1
XFILLER_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13250_ _13250_/A vssd1 vssd1 vccd1 vccd1 _14879_/A sky130_fd_sc_hd__buf_4
X_10462_ _10693_/A vssd1 vssd1 vccd1 vccd1 _10503_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ _15803_/Q _12369_/B _12208_/C vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__nand3_1
XFILLER_135_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _15959_/Q _13286_/B _13187_/C vssd1 vssd1 vccd1 vccd1 _13181_/Y sky130_fd_sc_hd__nand3_1
XFILLER_136_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10393_ _10391_/Y _10386_/C _10398_/A _10390_/Y vssd1 vssd1 vccd1 vccd1 _10398_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12132_ _12170_/A _12132_/B _12132_/C vssd1 vssd1 vccd1 vccd1 _12133_/A sky130_fd_sc_hd__and3_1
XFILLER_123_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12063_ _12631_/A vssd1 vssd1 vccd1 vccd1 _12063_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11014_ _15617_/Q _11244_/B _11021_/C vssd1 vssd1 vccd1 vccd1 _11014_/X sky130_fd_sc_hd__and3_1
XFILLER_77_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15822_ _15907_/CLK _15822_/D vssd1 vssd1 vccd1 vccd1 _15822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15753_ _15763_/CLK _15753_/D vssd1 vssd1 vccd1 vccd1 _15753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12965_ _12971_/A _12963_/Y _12964_/Y _12959_/C vssd1 vssd1 vccd1 vccd1 _12967_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11916_ _15758_/Q _12085_/B _11923_/C vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__nand3_1
X_14704_ _16256_/Q _14778_/B _14706_/C vssd1 vssd1 vccd1 vccd1 _14709_/A sky130_fd_sc_hd__and3_1
X_15684_ _15763_/CLK _15684_/D vssd1 vssd1 vccd1 vccd1 _15684_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12896_ _15912_/Q _14031_/A _12896_/C vssd1 vssd1 vccd1 vccd1 _12896_/Y sky130_fd_sc_hd__nand3_1
XFILLER_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14635_ hold23/A _14639_/C _07649_/X vssd1 vssd1 vccd1 vccd1 _14635_/Y sky130_fd_sc_hd__a21oi_1
X_11847_ _12418_/A vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _16223_/Q _14566_/B _14566_/C vssd1 vssd1 vccd1 vccd1 _14566_/X sky130_fd_sc_hd__and3_1
XFILLER_13_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11778_ _11778_/A _11778_/B vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__nor2_1
X_16305_ _16337_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 _16305_/Q sky130_fd_sc_hd__dfxtp_1
X_13517_ _13412_/X _13514_/C _13516_/Y vssd1 vssd1 vccd1 vccd1 _16016_/D sky130_fd_sc_hd__a21oi_1
X_10729_ _15571_/Q _10729_/B _10734_/C vssd1 vssd1 vccd1 vccd1 _10729_/Y sky130_fd_sc_hd__nand3_1
XFILLER_146_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14497_ _14325_/X _14493_/B _14326_/X vssd1 vssd1 vccd1 vccd1 _14499_/A sky130_fd_sc_hd__a21oi_1
XFILLER_146_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16236_ _16247_/CLK _16236_/D vssd1 vssd1 vccd1 vccd1 _16236_/Q sky130_fd_sc_hd__dfxtp_2
X_13448_ _13455_/A _13446_/Y _13447_/Y _13442_/C vssd1 vssd1 vccd1 vccd1 _13450_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16167_ _16169_/CLK _16167_/D vssd1 vssd1 vccd1 vccd1 _16167_/Q sky130_fd_sc_hd__dfxtp_1
X_13379_ _13379_/A vssd1 vssd1 vccd1 vccd1 _15992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15118_ _14964_/X _15120_/C _15086_/X vssd1 vssd1 vccd1 vccd1 _15119_/B sky130_fd_sc_hd__o21ai_1
XFILLER_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16098_ _16119_/CLK _16098_/D vssd1 vssd1 vccd1 vccd1 _16098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07940_ _08610_/C _07942_/B vssd1 vssd1 vccd1 vccd1 _08163_/A sky130_fd_sc_hd__nor2_2
X_15049_ _15049_/A _15049_/B vssd1 vssd1 vccd1 vccd1 _16329_/D sky130_fd_sc_hd__nor2_1
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07871_ _16071_/Q _16089_/Q vssd1 vssd1 vccd1 vccd1 _07873_/A sky130_fd_sc_hd__or2_1
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09610_ _15398_/Q _09615_/C _09490_/X vssd1 vssd1 vccd1 vccd1 _09612_/C sky130_fd_sc_hd__a21o_1
XFILLER_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09541_ _09541_/A vssd1 vssd1 vccd1 vccd1 _09541_/X sky130_fd_sc_hd__buf_2
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ _09472_/A _09476_/C vssd1 vssd1 vccd1 vccd1 _09472_/X sky130_fd_sc_hd__or2_1
XFILLER_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ state1[2] _08433_/A vssd1 vssd1 vccd1 vccd1 _08424_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08354_ _08295_/A _08295_/B _08353_/X vssd1 vssd1 vccd1 vccd1 _08356_/C sky130_fd_sc_hd__o21a_2
X_08285_ _08285_/A _08200_/A vssd1 vssd1 vccd1 vccd1 _08285_/X sky130_fd_sc_hd__or2b_1
XFILLER_117_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09808_ _09808_/A vssd1 vssd1 vccd1 vccd1 _15427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09739_ _09739_/A vssd1 vssd1 vccd1 vccd1 _15417_/D sky130_fd_sc_hd__clkbuf_1
X_12750_ _12757_/B _12750_/B vssd1 vssd1 vccd1 vccd1 _12752_/A sky130_fd_sc_hd__or2_1
XFILLER_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11701_/A vssd1 vssd1 vccd1 vccd1 _15723_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12681_/A vssd1 vssd1 vccd1 vccd1 _15877_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14420_/A _14420_/B vssd1 vssd1 vccd1 vccd1 _16187_/D sky130_fd_sc_hd__nor2_1
X_11632_ _11653_/A _11632_/B _11632_/C vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__and3_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14351_ _16177_/Q _14357_/C _14177_/X vssd1 vssd1 vccd1 vccd1 _14353_/B sky130_fd_sc_hd__a21oi_1
X_11563_ _11576_/C vssd1 vssd1 vccd1 vccd1 _11585_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13302_ _13457_/A _13304_/C vssd1 vssd1 vccd1 vccd1 _13302_/X sky130_fd_sc_hd__or2_1
X_10514_ _10520_/B _10514_/B vssd1 vssd1 vccd1 vccd1 _10516_/A sky130_fd_sc_hd__or2_1
XFILLER_10_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14282_ _14061_/X _14153_/X _14277_/B _14240_/X vssd1 vssd1 vccd1 vccd1 _14283_/B
+ sky130_fd_sc_hd__a31o_1
X_11494_ _11492_/A _11492_/B _11493_/X vssd1 vssd1 vccd1 vccd1 _15690_/D sky130_fd_sc_hd__a21oi_1
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16021_ _16031_/CLK _16021_/D vssd1 vssd1 vccd1 vccd1 _16021_/Q sky130_fd_sc_hd__dfxtp_1
X_13233_ _15969_/Q _13240_/C _13179_/X vssd1 vssd1 vccd1 vccd1 _13233_/Y sky130_fd_sc_hd__a21oi_1
X_10445_ _10445_/A vssd1 vssd1 vccd1 vccd1 _15526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ _13283_/A vssd1 vssd1 vccd1 vccd1 _13223_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _10372_/X _10374_/Y _10375_/Y _10368_/C vssd1 vssd1 vccd1 vccd1 _10378_/B
+ sky130_fd_sc_hd__o211ai_1
X_12115_ _15789_/Q _12228_/B _12115_/C vssd1 vssd1 vccd1 vccd1 _12124_/A sky130_fd_sc_hd__and3_1
X_13095_ _15948_/Q _13138_/C _13041_/X vssd1 vssd1 vccd1 vccd1 _13098_/B sky130_fd_sc_hd__a21oi_1
XFILLER_112_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12046_ _12046_/A vssd1 vssd1 vccd1 vccd1 _15777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _07603_/A _15805_/D vssd1 vssd1 vccd1 vccd1 _15805_/Q sky130_fd_sc_hd__dfxtp_1
X_13997_ _16105_/Q _14003_/C _13893_/X vssd1 vssd1 vccd1 vccd1 _13999_/B sky130_fd_sc_hd__a21oi_1
XFILLER_80_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15736_ _15763_/CLK _15736_/D vssd1 vssd1 vccd1 vccd1 _15736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12948_ _15922_/Q _12949_/C _13130_/A vssd1 vssd1 vccd1 vccd1 _12948_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15667_ _15763_/CLK _15667_/D vssd1 vssd1 vccd1 vccd1 _15667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12879_ _15910_/Q _12879_/B _12887_/C vssd1 vssd1 vccd1 vccd1 _12884_/A sky130_fd_sc_hd__and3_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14618_ _14368_/A _08541_/X _14612_/B _14459_/X vssd1 vssd1 vccd1 vccd1 _14619_/B
+ sky130_fd_sc_hd__a31o_1
X_15598_ _15194_/Q _15598_/D vssd1 vssd1 vccd1 vccd1 _15598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14549_ _16220_/Q _14554_/C _07632_/A vssd1 vssd1 vccd1 vccd1 _14551_/C sky130_fd_sc_hd__a21o_1
X_08070_ _15647_/Q vssd1 vssd1 vccd1 vccd1 _11213_/A sky130_fd_sc_hd__inv_2
XFILLER_146_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16219_ _16240_/CLK _16219_/D vssd1 vssd1 vccd1 vccd1 _16219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08972_ _09066_/A _08972_/B _08976_/A vssd1 vssd1 vccd1 vccd1 _15298_/D sky130_fd_sc_hd__nor3_1
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07923_ _10121_/A _07980_/B vssd1 vssd1 vccd1 vccd1 _07924_/B sky130_fd_sc_hd__xnor2_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07854_ _16125_/Q _16143_/Q vssd1 vssd1 vccd1 vccd1 _07996_/B sky130_fd_sc_hd__xor2_2
X_07785_ _11502_/A _07785_/B vssd1 vssd1 vccd1 vccd1 _07786_/B sky130_fd_sc_hd__xnor2_2
XFILLER_25_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09524_ _15383_/Q _09524_/B _09528_/C vssd1 vssd1 vccd1 vccd1 _09524_/Y sky130_fd_sc_hd__nand3_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09455_ _15373_/Q _09572_/B _09460_/C vssd1 vssd1 vccd1 vccd1 _09455_/Y sky130_fd_sc_hd__nand3_1
XFILLER_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08406_ _08389_/A _08389_/B _08387_/A vssd1 vssd1 vccd1 vccd1 _08406_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09386_ _15364_/Q _09444_/B _09391_/C vssd1 vssd1 vccd1 vccd1 _09386_/X sky130_fd_sc_hd__and3_1
X_08337_ _08331_/Y _08333_/X _08336_/Y vssd1 vssd1 vccd1 vccd1 _15209_/D sky130_fd_sc_hd__a21oi_1
XFILLER_137_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08268_ _08268_/A _08282_/A vssd1 vssd1 vccd1 vccd1 _08270_/C sky130_fd_sc_hd__xor2_4
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08199_ _08199_/A _08199_/B vssd1 vssd1 vccd1 vccd1 _08285_/A sky130_fd_sc_hd__xnor2_2
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10230_ _10266_/A _10230_/B _10230_/C vssd1 vssd1 vccd1 vccd1 _10231_/A sky130_fd_sc_hd__and3_1
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10161_ _10219_/A _10161_/B _10165_/B vssd1 vssd1 vccd1 vccd1 _15482_/D sky130_fd_sc_hd__nor3_1
XFILLER_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _15473_/Q _10317_/B _10100_/C vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__and3_1
XFILLER_102_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13920_ _13920_/A vssd1 vssd1 vccd1 vccd1 _13920_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13851_ _13849_/Y _13844_/C _13856_/A _13848_/Y vssd1 vssd1 vccd1 vccd1 _13856_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12802_ _12808_/A _12799_/Y _12801_/Y _12796_/C vssd1 vssd1 vccd1 vccd1 _12804_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13782_ _13782_/A _13782_/B _13782_/C vssd1 vssd1 vccd1 vccd1 _13783_/C sky130_fd_sc_hd__nand3_1
XFILLER_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10994_ _15614_/Q _10999_/C _10933_/X vssd1 vssd1 vccd1 vccd1 _10996_/C sky130_fd_sc_hd__a21o_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15521_ _15539_/CLK _15521_/D vssd1 vssd1 vccd1 vccd1 _15521_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _12733_/A vssd1 vssd1 vccd1 vccd1 _15885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _15483_/CLK _15452_/D vssd1 vssd1 vccd1 vccd1 _15452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12657_/B _12658_/C _12660_/X _12662_/Y vssd1 vssd1 vccd1 vccd1 _12665_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _16187_/Q _14566_/B _14403_/C vssd1 vssd1 vccd1 vccd1 _14403_/X sky130_fd_sc_hd__and3_1
X_11615_ _12188_/A vssd1 vssd1 vccd1 vccd1 _11615_/X sky130_fd_sc_hd__clkbuf_2
X_15383_ _15484_/CLK _15383_/D vssd1 vssd1 vccd1 vccd1 _15383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12595_ _15866_/Q _12653_/B _12601_/C vssd1 vssd1 vccd1 vccd1 _12598_/B sky130_fd_sc_hd__nand3_1
XFILLER_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14334_ _14337_/C vssd1 vssd1 vccd1 vccd1 _14345_/C sky130_fd_sc_hd__clkbuf_1
X_11546_ _11661_/A _11546_/B _11550_/B vssd1 vssd1 vccd1 vccd1 _15698_/D sky130_fd_sc_hd__nor3_1
XFILLER_51_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14265_ _14265_/A _14265_/B vssd1 vssd1 vccd1 vccd1 _14265_/X sky130_fd_sc_hd__or2_1
XFILLER_7_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11477_ _11477_/A _11477_/B _11477_/C vssd1 vssd1 vccd1 vccd1 _11478_/A sky130_fd_sc_hd__and3_1
XFILLER_109_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16004_ _16011_/CLK _16004_/D vssd1 vssd1 vccd1 vccd1 _16004_/Q sky130_fd_sc_hd__dfxtp_1
X_13216_ _13474_/A vssd1 vssd1 vccd1 vccd1 _13420_/B sky130_fd_sc_hd__buf_2
X_10428_ _10426_/X _10427_/Y _10421_/B _10422_/C vssd1 vssd1 vccd1 vccd1 _10430_/B
+ sky130_fd_sc_hd__o211ai_1
X_14196_ _14316_/A vssd1 vssd1 vccd1 vccd1 _14196_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13147_ _14653_/A vssd1 vssd1 vccd1 vccd1 _14892_/A sky130_fd_sc_hd__buf_4
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _10360_/B _10360_/C _10360_/A vssd1 vssd1 vccd1 vccd1 _10361_/B sky130_fd_sc_hd__a21o_1
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _15944_/Q _13078_/B _13078_/C vssd1 vssd1 vccd1 vccd1 _13086_/B sky130_fd_sc_hd__and3_1
XFILLER_111_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12029_ _12030_/B _12030_/C _12030_/A vssd1 vssd1 vccd1 vccd1 _12031_/B sky130_fd_sc_hd__a21o_1
XFILLER_78_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15719_ _15728_/CLK _15719_/D vssd1 vssd1 vccd1 vccd1 _15719_/Q sky130_fd_sc_hd__dfxtp_1
X_09240_ _09238_/Y _09233_/C _09245_/A _09237_/Y vssd1 vssd1 vccd1 vccd1 _09245_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ _09171_/A _09171_/B _09171_/C vssd1 vssd1 vccd1 vccd1 _09172_/A sky130_fd_sc_hd__and3_1
XFILLER_119_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08122_ _08242_/A _08242_/B vssd1 vssd1 vccd1 vccd1 _08131_/A sky130_fd_sc_hd__xor2_4
XFILLER_119_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ _08211_/A _08053_/B vssd1 vssd1 vccd1 vccd1 _08064_/A sky130_fd_sc_hd__and2_2
XFILLER_127_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08955_ _13930_/A vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07906_ _16269_/Q _07963_/A _07906_/C vssd1 vssd1 vccd1 vccd1 _07963_/B sky130_fd_sc_hd__nand3_4
X_08886_ _15287_/Q _09067_/B _08886_/C vssd1 vssd1 vccd1 vccd1 _08897_/B sky130_fd_sc_hd__and3_1
X_07837_ _15899_/Q _08030_/B vssd1 vssd1 vccd1 vccd1 _08025_/B sky130_fd_sc_hd__xnor2_2
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07768_ _15611_/Q _15593_/Q vssd1 vssd1 vccd1 vccd1 _07771_/B sky130_fd_sc_hd__or2_1
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _15382_/Q _09508_/C _09506_/X vssd1 vssd1 vccd1 vccd1 _09507_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _13715_/A vssd1 vssd1 vccd1 vccd1 _14653_/A sky130_fd_sc_hd__buf_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _15372_/Q _09496_/B _09438_/C vssd1 vssd1 vccd1 vccd1 _09438_/X sky130_fd_sc_hd__and3_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _09391_/C vssd1 vssd1 vccd1 vccd1 _09403_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11400_ _11400_/A vssd1 vssd1 vccd1 vccd1 _15676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12380_ _12373_/B _12374_/C _12376_/X _12378_/Y vssd1 vssd1 vccd1 vccd1 _12381_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11331_ _15673_/Q _15672_/Q _15671_/Q _11273_/X vssd1 vssd1 vccd1 vccd1 _15665_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_119_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14050_ _14045_/Y _14048_/X _14049_/X vssd1 vssd1 vccd1 vccd1 _14050_/Y sky130_fd_sc_hd__a21oi_1
X_11262_ _11262_/A _11262_/B vssd1 vssd1 vccd1 vccd1 _11264_/B sky130_fd_sc_hd__nor2_1
X_13001_ _13001_/A vssd1 vssd1 vccd1 vccd1 _15929_/D sky130_fd_sc_hd__clkbuf_1
X_10213_ _11422_/A vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_97_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11193_ _15644_/Q _11313_/B _11198_/C vssd1 vssd1 vccd1 vccd1 _11193_/Y sky130_fd_sc_hd__nand3_1
X_10144_ _10141_/X _10142_/Y _10143_/Y _10139_/C vssd1 vssd1 vccd1 vccd1 _10146_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10075_ _10940_/A vssd1 vssd1 vccd1 vccd1 _10075_/X sky130_fd_sc_hd__clkbuf_2
X_14952_ _15023_/A _14952_/B _14956_/B vssd1 vssd1 vccd1 vccd1 _16308_/D sky130_fd_sc_hd__nor3_1
XFILLER_121_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13903_ _16088_/Q _14137_/B _13903_/C vssd1 vssd1 vccd1 vccd1 _13903_/X sky130_fd_sc_hd__and3_1
X_14883_ _14883_/A vssd1 vssd1 vccd1 vccd1 _15045_/A sky130_fd_sc_hd__buf_2
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13834_ _13832_/X _13833_/Y _13829_/B _13830_/C vssd1 vssd1 vccd1 vccd1 _13836_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _13763_/A _13763_/B _13764_/X vssd1 vssd1 vccd1 vccd1 _16059_/D sky130_fd_sc_hd__a21oi_1
X_10977_ _10975_/A _10975_/B _10976_/X vssd1 vssd1 vccd1 vccd1 _15609_/D sky130_fd_sc_hd__a21oi_1
X_15504_ _15224_/Q _15504_/D vssd1 vssd1 vccd1 vccd1 _15504_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12716_ _12717_/B _12717_/C _12717_/A vssd1 vssd1 vccd1 vccd1 _12718_/B sky130_fd_sc_hd__a21o_1
X_13696_ _13692_/X _13694_/Y _13695_/Y _13690_/C vssd1 vssd1 vccd1 vccd1 _13698_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15435_ _15483_/CLK _15435_/D vssd1 vssd1 vccd1 vccd1 _15435_/Q sky130_fd_sc_hd__dfxtp_1
X_12647_ _12670_/C vssd1 vssd1 vccd1 vccd1 _12684_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15366_ _15440_/CLK _15366_/D vssd1 vssd1 vccd1 vccd1 _15366_/Q sky130_fd_sc_hd__dfxtp_1
X_12578_ _12578_/A _12578_/B vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14317_ _14312_/Y _14315_/X _14316_/X vssd1 vssd1 vccd1 vccd1 _14317_/Y sky130_fd_sc_hd__a21oi_1
X_11529_ _11525_/X _11527_/Y _11528_/Y _11523_/C vssd1 vssd1 vccd1 vccd1 _11531_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15297_ _15449_/CLK _15297_/D vssd1 vssd1 vccd1 vccd1 _15297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14248_ _14304_/A _14248_/B _14253_/A vssd1 vssd1 vccd1 vccd1 _16153_/D sky130_fd_sc_hd__nor3_1
X_14179_ _14179_/A _14179_/B vssd1 vssd1 vccd1 vccd1 _14179_/Y sky130_fd_sc_hd__nor2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _15264_/Q _08745_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _08742_/C sky130_fd_sc_hd__a21o_1
XFILLER_79_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08671_ _15269_/Q _15268_/Q _15267_/Q _08604_/X vssd1 vssd1 vccd1 vccd1 _15252_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_94_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07622_ _14901_/A vssd1 vssd1 vccd1 vccd1 _08735_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09223_ _09219_/X _09221_/Y _09222_/Y _09216_/C vssd1 vssd1 vccd1 vccd1 _09225_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_139_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09154_ _09152_/X _09153_/Y _09149_/B _09150_/C vssd1 vssd1 vccd1 vccd1 _09156_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08105_ _08105_/A _08225_/A vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__xnor2_4
X_09085_ _09105_/C vssd1 vssd1 vccd1 vccd1 _09117_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08036_ _08214_/B _08036_/B vssd1 vssd1 vccd1 vccd1 _08037_/B sky130_fd_sc_hd__xnor2_2
XFILLER_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09987_ input7/X vssd1 vssd1 vccd1 vccd1 _11197_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08938_ _15294_/Q _08945_/C _08873_/X vssd1 vssd1 vccd1 vccd1 _08938_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08869_ _08867_/Y _08863_/C _08865_/X _08866_/Y vssd1 vssd1 vccd1 vccd1 _08870_/C
+ sky130_fd_sc_hd__a211o_1
X_10900_ _10895_/X _10898_/Y _10899_/Y _10893_/C vssd1 vssd1 vccd1 vccd1 _10902_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_45_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11880_ _15751_/Q _11938_/B _11885_/C vssd1 vssd1 vccd1 vccd1 _11880_/Y sky130_fd_sc_hd__nand3_1
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10831_ _15589_/Q _10888_/B _10835_/C vssd1 vssd1 vccd1 vccd1 _10831_/X sky130_fd_sc_hd__and3_1
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ _16023_/Q _13550_/B _13554_/C vssd1 vssd1 vccd1 vccd1 _13550_/Y sky130_fd_sc_hd__nand3_1
Xrepeater16 _15224_/Q vssd1 vssd1 vccd1 vccd1 _15484_/CLK sky130_fd_sc_hd__buf_12
X_10762_ _15577_/Q _10817_/B _10770_/C vssd1 vssd1 vccd1 vccd1 _10767_/A sky130_fd_sc_hd__and3_1
X_12501_ _12498_/X _12499_/Y _12500_/Y _12496_/C vssd1 vssd1 vccd1 vccd1 _12503_/B
+ sky130_fd_sc_hd__o211ai_1
X_13481_ _13481_/A _13481_/B _13481_/C vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__and3_1
X_10693_ _10693_/A vssd1 vssd1 vccd1 vccd1 _10732_/A sky130_fd_sc_hd__clkbuf_2
X_15220_ _16242_/CLK _15220_/D vssd1 vssd1 vccd1 vccd1 state1[5] sky130_fd_sc_hd__dfxtp_2
X_12432_ _12454_/A _12432_/B _12432_/C vssd1 vssd1 vccd1 vccd1 _12433_/A sky130_fd_sc_hd__and3_1
XFILLER_139_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15151_ _15001_/X _15144_/A _15147_/B _15150_/Y vssd1 vssd1 vccd1 vccd1 _16355_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _12386_/C vssd1 vssd1 vccd1 vccd1 _12399_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _14102_/A _14102_/B vssd1 vssd1 vccd1 vccd1 _14103_/B sky130_fd_sc_hd__nor2_1
X_11314_ _11320_/A _11312_/Y _11313_/Y _11309_/C vssd1 vssd1 vccd1 vccd1 _11316_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15082_ _15152_/A _15085_/C vssd1 vssd1 vccd1 vccd1 _15084_/A sky130_fd_sc_hd__and2_1
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12294_ _12294_/A _12294_/B vssd1 vssd1 vccd1 vccd1 _12295_/B sky130_fd_sc_hd__nor2_1
XFILLER_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14033_ _14300_/A vssd1 vssd1 vccd1 vccd1 _14033_/X sky130_fd_sc_hd__clkbuf_2
X_11245_ _15653_/Q _11253_/C _11184_/X vssd1 vssd1 vccd1 vccd1 _11245_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _15643_/Q _11178_/C _10948_/X vssd1 vssd1 vccd1 vccd1 _11176_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10127_ _10219_/A _10127_/B _10131_/A vssd1 vssd1 vccd1 vccd1 _15477_/D sky130_fd_sc_hd__nor3_1
X_15984_ _15984_/CLK _15984_/D vssd1 vssd1 vccd1 vccd1 _15984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10058_ _10058_/A vssd1 vssd1 vccd1 vccd1 _10074_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14935_ hold6/X hold5/X _16320_/Q _14818_/X vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__o31a_1
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14866_ _14866_/A _14866_/B _14866_/C vssd1 vssd1 vccd1 vccd1 _14867_/C sky130_fd_sc_hd__nand3_1
XFILLER_91_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13817_ _13666_/X _13814_/C _13816_/Y vssd1 vssd1 vccd1 vccd1 _16070_/D sky130_fd_sc_hd__a21oi_1
XFILLER_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14797_ _14797_/A _14797_/B vssd1 vssd1 vccd1 vccd1 _14799_/A sky130_fd_sc_hd__or2_1
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13748_ _13746_/Y _13742_/C _13744_/X _13745_/Y vssd1 vssd1 vccd1 vccd1 _13749_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13679_ _13679_/A vssd1 vssd1 vccd1 vccd1 _14074_/B sky130_fd_sc_hd__buf_2
X_15418_ _15483_/CLK _15418_/D vssd1 vssd1 vccd1 vccd1 _15418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15349_ _15368_/CLK _15349_/D vssd1 vssd1 vccd1 vccd1 _15349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09910_ _15445_/Q _09911_/C _09794_/X vssd1 vssd1 vccd1 vccd1 _09910_/Y sky130_fd_sc_hd__a21oi_1
X_09841_ _15434_/Q _09847_/C _09778_/X vssd1 vssd1 vccd1 vccd1 _09843_/C sky130_fd_sc_hd__a21o_1
XFILLER_98_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09811_/C vssd1 vssd1 vccd1 vccd1 _09817_/C sky130_fd_sc_hd__clkbuf_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08765_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08654_ _08660_/A _08652_/Y _08653_/Y _08648_/C vssd1 vssd1 vccd1 vccd1 _08656_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ _11898_/A vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__buf_2
X_08585_ _08593_/A _08583_/Y _08584_/Y _08580_/C vssd1 vssd1 vccd1 vccd1 _08587_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09206_ _15336_/Q _09211_/C _09205_/X vssd1 vssd1 vccd1 vccd1 _09208_/C sky130_fd_sc_hd__a21o_1
X_09137_ _15341_/Q _15340_/Q _15339_/Q _08901_/X vssd1 vssd1 vccd1 vccd1 _15324_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_135_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _15314_/Q _09067_/C _08888_/X vssd1 vssd1 vccd1 vccd1 _09069_/B sky130_fd_sc_hd__a21oi_1
XFILLER_135_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08019_ _08019_/A _08019_/B vssd1 vssd1 vccd1 vccd1 _08020_/B sky130_fd_sc_hd__and2_1
XFILLER_135_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11030_ _11030_/A _11030_/B vssd1 vssd1 vccd1 vccd1 _11031_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12981_ _13723_/A vssd1 vssd1 vccd1 vccd1 _12981_/X sky130_fd_sc_hd__buf_2
X_14720_ _14720_/A _14720_/B vssd1 vssd1 vccd1 vccd1 _14722_/A sky130_fd_sc_hd__or2_1
X_11932_ _11929_/X _11930_/Y _11931_/Y _11927_/C vssd1 vssd1 vccd1 vccd1 _11934_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11863_ _15750_/Q _11863_/B _11863_/C vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__and3_1
X_14651_ _07688_/X _14654_/C _07690_/X vssd1 vssd1 vccd1 vccd1 _14652_/B sky130_fd_sc_hd__o21ai_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10814_ _10835_/C vssd1 vssd1 vccd1 vccd1 _10847_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13602_ _13608_/A _13599_/Y _13601_/Y _13595_/C vssd1 vssd1 vccd1 vccd1 _13604_/B
+ sky130_fd_sc_hd__o211a_1
X_11794_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12025_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14582_ _14593_/C vssd1 vssd1 vccd1 vccd1 _14605_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16321_ _16321_/CLK _16321_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
X_13533_ _16022_/Q _13738_/B _13533_/C vssd1 vssd1 vccd1 vccd1 _13533_/X sky130_fd_sc_hd__and3_1
X_10745_ _10745_/A _10745_/B vssd1 vssd1 vccd1 vccd1 _10750_/C sky130_fd_sc_hd__nor2_1
XFILLER_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13464_ _15086_/A vssd1 vssd1 vccd1 vccd1 _13464_/X sky130_fd_sc_hd__clkbuf_2
X_16252_ _16264_/CLK _16252_/D vssd1 vssd1 vccd1 vccd1 _16252_/Q sky130_fd_sc_hd__dfxtp_2
X_10676_ _10676_/A _10676_/B _10676_/C vssd1 vssd1 vccd1 vccd1 _10677_/A sky130_fd_sc_hd__and3_1
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12415_ _12414_/B _12414_/C _12188_/X vssd1 vssd1 vccd1 vccd1 _12416_/C sky130_fd_sc_hd__o21ai_1
X_15203_ _16241_/CLK _15203_/D vssd1 vssd1 vccd1 vccd1 _15203_/Q sky130_fd_sc_hd__dfxtp_1
X_16183_ _16192_/CLK _16183_/D vssd1 vssd1 vccd1 vccd1 _16183_/Q sky130_fd_sc_hd__dfxtp_1
X_13395_ _15997_/Q _13401_/C _13342_/X vssd1 vssd1 vccd1 vccd1 _13395_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15134_ _15134_/A _15134_/B _15134_/C vssd1 vssd1 vccd1 vccd1 _15135_/C sky130_fd_sc_hd__nand3_1
X_12346_ _15826_/Q _12575_/B _12346_/C vssd1 vssd1 vccd1 vccd1 _12356_/B sky130_fd_sc_hd__and3_1
XFILLER_142_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15065_ _15135_/A _15065_/B _15065_/C vssd1 vssd1 vccd1 vccd1 _15066_/A sky130_fd_sc_hd__and3_1
X_12277_ _12277_/A vssd1 vssd1 vccd1 vccd1 _12507_/B sky130_fd_sc_hd__buf_2
XFILLER_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14016_ _14413_/A _15013_/A _14011_/B _13969_/X vssd1 vssd1 vccd1 vccd1 _14017_/B
+ sky130_fd_sc_hd__a31o_1
X_11228_ _15651_/Q _11289_/B _11228_/C vssd1 vssd1 vccd1 vccd1 _11228_/X sky130_fd_sc_hd__and3_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11159_ _11191_/C vssd1 vssd1 vccd1 vccd1 _11198_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15967_ _16123_/CLK _15967_/D vssd1 vssd1 vccd1 vccd1 _15967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14918_ hold17/X _14916_/C _14917_/X vssd1 vssd1 vccd1 vccd1 _14919_/B sky130_fd_sc_hd__a21oi_1
X_15898_ _07603_/A _15898_/D vssd1 vssd1 vccd1 vccd1 _15898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14849_ _14963_/A _14853_/C vssd1 vssd1 vccd1 vccd1 _14851_/A sky130_fd_sc_hd__and2_1
XFILLER_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _08442_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08372_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09824_ _09822_/A _09822_/B _09823_/X vssd1 vssd1 vccd1 vccd1 _15429_/D sky130_fd_sc_hd__a21oi_1
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09755_ _10044_/A vssd1 vssd1 vccd1 vccd1 _09755_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08706_ _15259_/Q _10963_/C _08706_/C vssd1 vssd1 vccd1 vccd1 _08718_/A sky130_fd_sc_hd__and3_1
X_09686_ _15410_/Q _09692_/C _09453_/X vssd1 vssd1 vccd1 vccd1 _09686_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _08632_/X _08635_/Y _08636_/Y _08629_/C vssd1 vssd1 vccd1 vccd1 _08639_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08568_ _15238_/Q _08753_/B _08568_/C vssd1 vssd1 vccd1 vccd1 _08568_/Y sky130_fd_sc_hd__nand3_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08499_ _10947_/A vssd1 vssd1 vccd1 vccd1 _11128_/A sky130_fd_sc_hd__buf_2
X_10530_ _10561_/C vssd1 vssd1 vccd1 vccd1 _10569_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_109_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _11612_/A vssd1 vssd1 vccd1 vccd1 _10693_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12200_ _12234_/A _12200_/B _12204_/A vssd1 vssd1 vccd1 vccd1 _15801_/D sky130_fd_sc_hd__nor3_1
XFILLER_108_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ _15960_/Q _13187_/C _13179_/X vssd1 vssd1 vccd1 vccd1 _13180_/Y sky130_fd_sc_hd__a21oi_1
X_10392_ _10398_/A _10390_/Y _10391_/Y _10386_/C vssd1 vssd1 vccd1 vccd1 _10394_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12131_ _12130_/B _12130_/C _11902_/X vssd1 vssd1 vccd1 vccd1 _12132_/C sky130_fd_sc_hd__o21ai_1
XFILLER_124_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ _15781_/Q _12291_/B _12062_/C vssd1 vssd1 vccd1 vccd1 _12072_/B sky130_fd_sc_hd__and3_1
XFILLER_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11013_ _11303_/A vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15821_ _07603_/A _15821_/D vssd1 vssd1 vccd1 vccd1 _15821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15752_ _15763_/CLK _15752_/D vssd1 vssd1 vccd1 vccd1 _15752_/Q sky130_fd_sc_hd__dfxtp_1
X_12964_ _15923_/Q _13018_/B _12968_/C vssd1 vssd1 vccd1 vccd1 _12964_/Y sky130_fd_sc_hd__nand3_1
XFILLER_45_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14703_ _16256_/Q _14717_/C _14702_/X vssd1 vssd1 vccd1 vccd1 _14705_/B sky130_fd_sc_hd__a21oi_1
X_11915_ _11949_/A _11915_/B _11919_/A vssd1 vssd1 vccd1 vccd1 _15756_/D sky130_fd_sc_hd__nor3_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15683_/CLK _15683_/D vssd1 vssd1 vccd1 vccd1 _15683_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12895_ _13532_/A vssd1 vssd1 vccd1 vccd1 _14031_/A sky130_fd_sc_hd__buf_4
XFILLER_60_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14634_ hold23/A _14634_/B _14639_/C vssd1 vssd1 vccd1 vccd1 _14642_/A sky130_fd_sc_hd__and3_1
X_11846_ _11846_/A vssd1 vssd1 vccd1 vccd1 _15745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11777_ _11784_/B _11777_/B vssd1 vssd1 vccd1 vccd1 _11779_/A sky130_fd_sc_hd__or2_1
X_14565_ _14562_/B _14561_/Y _14562_/A vssd1 vssd1 vccd1 vccd1 _14565_/Y sky130_fd_sc_hd__o21bai_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16304_ _16304_/CLK _16304_/D vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
X_10728_ _15572_/Q _10734_/C _10610_/X vssd1 vssd1 vccd1 vccd1 _10728_/Y sky130_fd_sc_hd__a21oi_1
X_13516_ _13362_/X _13514_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13516_/Y sky130_fd_sc_hd__o21ai_1
X_14496_ _14413_/X _14493_/B _14495_/Y vssd1 vssd1 vccd1 vccd1 _16204_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16235_ _16247_/CLK _16235_/D vssd1 vssd1 vccd1 vccd1 _16235_/Q sky130_fd_sc_hd__dfxtp_2
X_10659_ _10676_/A _10659_/B _10659_/C vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__and3_1
XFILLER_127_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13447_ _16005_/Q _13550_/B _13451_/C vssd1 vssd1 vccd1 vccd1 _13447_/Y sky130_fd_sc_hd__nand3_1
XFILLER_70_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16166_ _16166_/CLK _16166_/D vssd1 vssd1 vccd1 vccd1 _16166_/Q sky130_fd_sc_hd__dfxtp_1
X_13378_ _13410_/A _13378_/B _13378_/C vssd1 vssd1 vccd1 vccd1 _13379_/A sky130_fd_sc_hd__and3_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15117_ _15152_/A _15120_/C vssd1 vssd1 vccd1 vccd1 _15119_/A sky130_fd_sc_hd__and2_1
X_12329_ _12337_/A _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _12330_/A sky130_fd_sc_hd__and3_1
X_16097_ _16367_/CLK _16097_/D vssd1 vssd1 vccd1 vccd1 _16097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15048_ _14964_/X _15051_/C _15007_/X vssd1 vssd1 vccd1 vccd1 _15049_/B sky130_fd_sc_hd__o21ai_1
X_07870_ _16107_/Q vssd1 vssd1 vccd1 vccd1 _14584_/C sky130_fd_sc_hd__inv_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09540_ _09540_/A vssd1 vssd1 vccd1 vccd1 _15385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09471_ _09471_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09476_/C sky130_fd_sc_hd__nor2_1
XFILLER_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08422_ spike_out[0] vssd1 vssd1 vccd1 vccd1 _08433_/A sky130_fd_sc_hd__inv_2
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08353_ _08293_/A _08293_/B _08296_/B vssd1 vssd1 vccd1 vccd1 _08353_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08284_ _08266_/A _08266_/B _08283_/X vssd1 vssd1 vccd1 vccd1 _08338_/B sky130_fd_sc_hd__o21ai_4
XFILLER_20_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09807_ _09807_/A _09807_/B _09807_/C vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__and3_1
XFILLER_75_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07999_ _07999_/A _07999_/B vssd1 vssd1 vccd1 vccd1 _08000_/B sky130_fd_sc_hd__or2_1
XFILLER_28_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09738_ _09746_/A _09738_/B _09738_/C vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__and3_1
XFILLER_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09669_ _09690_/A _09669_/B _09669_/C vssd1 vssd1 vccd1 vccd1 _09670_/A sky130_fd_sc_hd__and3_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11708_/A _11700_/B _11700_/C vssd1 vssd1 vccd1 vccd1 _11701_/A sky130_fd_sc_hd__and3_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12680_ _12680_/A _12680_/B _12680_/C vssd1 vssd1 vccd1 vccd1 _12681_/A sky130_fd_sc_hd__and3_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11631_/A _11631_/B _11631_/C vssd1 vssd1 vccd1 vccd1 _11632_/C sky130_fd_sc_hd__nand3_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14350_ _16177_/Q _14440_/B _14357_/C vssd1 vssd1 vccd1 vccd1 _14353_/A sky130_fd_sc_hd__and3_1
X_11562_ _11562_/A vssd1 vssd1 vccd1 vccd1 _11576_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ _15538_/Q _10512_/C _10333_/X vssd1 vssd1 vccd1 vccd1 _10514_/B sky130_fd_sc_hd__a21oi_1
X_13301_ _13301_/A _13301_/B vssd1 vssd1 vccd1 vccd1 _13304_/C sky130_fd_sc_hd__nor2_1
X_14281_ _14058_/X _14277_/B _14059_/X vssd1 vssd1 vccd1 vccd1 _14283_/A sky130_fd_sc_hd__a21oi_1
X_11493_ _11493_/A _11497_/C vssd1 vssd1 vccd1 vccd1 _11493_/X sky130_fd_sc_hd__or2_1
XFILLER_109_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13232_ _15969_/Q _13333_/B _13240_/C vssd1 vssd1 vccd1 vccd1 _13232_/X sky130_fd_sc_hd__and3_1
X_16020_ _16031_/CLK _16020_/D vssd1 vssd1 vccd1 vccd1 _16020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10444_ _10444_/A _10444_/B _10444_/C vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__and3_1
XFILLER_136_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ _13218_/A _13163_/B _13169_/A vssd1 vssd1 vccd1 vccd1 _15955_/D sky130_fd_sc_hd__nor3_1
XFILLER_123_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10375_ _15516_/Q _10492_/B _10375_/C vssd1 vssd1 vccd1 vccd1 _10375_/Y sky130_fd_sc_hd__nand3_1
X_12114_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__buf_2
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13094_ _13127_/C vssd1 vssd1 vccd1 vccd1 _13138_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12045_ _12053_/A _12045_/B _12045_/C vssd1 vssd1 vccd1 vccd1 _12046_/A sky130_fd_sc_hd__and3_1
XFILLER_78_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15804_ _07603_/A _15804_/D vssd1 vssd1 vccd1 vccd1 _15804_/Q sky130_fd_sc_hd__dfxtp_1
X_13996_ _16105_/Q _14221_/B _14003_/C vssd1 vssd1 vccd1 vccd1 _13999_/A sky130_fd_sc_hd__and3_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15735_ _15763_/CLK _15735_/D vssd1 vssd1 vccd1 vccd1 _15735_/Q sky130_fd_sc_hd__dfxtp_1
X_12947_ _15922_/Q _12947_/B _12949_/C vssd1 vssd1 vccd1 vccd1 _12947_/X sky130_fd_sc_hd__and3_1
XFILLER_34_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15666_ _15763_/CLK _15666_/D vssd1 vssd1 vccd1 vccd1 _15666_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _15910_/Q _12914_/C _12767_/X vssd1 vssd1 vccd1 vccd1 _12880_/B sky130_fd_sc_hd__a21oi_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _07701_/X _14612_/B _14814_/A vssd1 vssd1 vccd1 vccd1 _14619_/A sky130_fd_sc_hd__a21oi_1
X_11829_ _15743_/Q _11887_/B _11833_/C vssd1 vssd1 vccd1 vccd1 _11829_/Y sky130_fd_sc_hd__nand3_1
X_15597_ _15194_/Q _15597_/D vssd1 vssd1 vccd1 vccd1 _15597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14548_ _16220_/Q _14587_/B _14554_/C vssd1 vssd1 vccd1 vccd1 _14551_/B sky130_fd_sc_hd__nand3_1
XFILLER_146_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14479_ _16204_/Q _14598_/B _14486_/C vssd1 vssd1 vccd1 vccd1 _14482_/A sky130_fd_sc_hd__and3_1
X_16218_ _16241_/CLK _16218_/D vssd1 vssd1 vccd1 vccd1 _16218_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_114_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16149_ _16169_/CLK _16149_/D vssd1 vssd1 vccd1 vccd1 _16149_/Q sky130_fd_sc_hd__dfxtp_1
X_08971_ _15299_/Q _09088_/B _08981_/C vssd1 vssd1 vccd1 vccd1 _08976_/A sky130_fd_sc_hd__and3_1
X_07922_ _10812_/A _07922_/B vssd1 vssd1 vccd1 vccd1 _07980_/B sky130_fd_sc_hd__xnor2_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07853_ _16062_/Q vssd1 vssd1 vccd1 vccd1 _13824_/C sky130_fd_sc_hd__clkinv_2
XFILLER_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07784_ _07784_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _07785_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09523_ _15384_/Q _09528_/C _09404_/X vssd1 vssd1 vccd1 vccd1 _09523_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09454_ _15374_/Q _09460_/C _09453_/X vssd1 vssd1 vccd1 vccd1 _09454_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08405_ _08393_/A _08393_/B _08404_/X vssd1 vssd1 vccd1 vccd1 _08414_/A sky130_fd_sc_hd__a21oi_2
X_09385_ _09385_/A vssd1 vssd1 vccd1 vccd1 _15362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08336_ _08331_/Y _08333_/X _08335_/X vssd1 vssd1 vccd1 vccd1 _08336_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08267_ _08267_/A _08283_/A vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__xor2_4
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08198_ _08198_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08199_/B sky130_fd_sc_hd__xor2_2
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10160_ _10158_/Y _10153_/C _10165_/A _10156_/Y vssd1 vssd1 vccd1 vccd1 _10165_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10091_ _11303_/A vssd1 vssd1 vccd1 vccd1 _10317_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13850_ _13856_/A _13848_/Y _13849_/Y _13844_/C vssd1 vssd1 vccd1 vccd1 _13852_/B
+ sky130_fd_sc_hd__o211a_1
X_12801_ _15896_/Q _13018_/B _12805_/C vssd1 vssd1 vccd1 vccd1 _12801_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13781_ _13782_/B _13782_/C _13782_/A vssd1 vssd1 vccd1 vccd1 _13783_/B sky130_fd_sc_hd__a21o_1
XFILLER_28_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10993_ _15614_/Q _11221_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _10996_/B sky130_fd_sc_hd__nand3_1
XFILLER_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15520_ _15655_/CLK _15520_/D vssd1 vssd1 vccd1 vccd1 _15520_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12740_/A _12732_/B _12732_/C vssd1 vssd1 vccd1 vccd1 _12733_/A sky130_fd_sc_hd__and3_1
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15451_ _15483_/CLK _15451_/D vssd1 vssd1 vccd1 vccd1 _15451_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12660_/X _12662_/Y _12657_/B _12658_/C vssd1 vssd1 vccd1 vccd1 _12665_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _14402_/A vssd1 vssd1 vccd1 vccd1 _14566_/B sky130_fd_sc_hd__clkbuf_2
X_11614_ _11727_/A _11614_/B _11614_/C vssd1 vssd1 vccd1 vccd1 _11617_/B sky130_fd_sc_hd__or3_1
X_15382_ _15484_/CLK _15382_/D vssd1 vssd1 vccd1 vccd1 _15382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12652_/A _12594_/B _12598_/A vssd1 vssd1 vccd1 vccd1 _15864_/D sky130_fd_sc_hd__nor3_1
X_14333_ _16161_/Q vssd1 vssd1 vccd1 vccd1 _14337_/C sky130_fd_sc_hd__inv_2
XFILLER_128_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11545_ _11543_/Y _11538_/C _11550_/A _11542_/Y vssd1 vssd1 vccd1 vccd1 _11550_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_11_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14264_ _14264_/A _14264_/B vssd1 vssd1 vccd1 vccd1 _14264_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11476_ _11474_/Y _11469_/C _11471_/X _11473_/Y vssd1 vssd1 vccd1 vccd1 _11477_/C
+ sky130_fd_sc_hd__a211o_1
X_16003_ _16011_/CLK _16003_/D vssd1 vssd1 vccd1 vccd1 _16003_/Q sky130_fd_sc_hd__dfxtp_1
X_10427_ _15525_/Q _10434_/C _10364_/X vssd1 vssd1 vccd1 vccd1 _10427_/Y sky130_fd_sc_hd__a21oi_1
X_13215_ _15966_/Q _13246_/C _13041_/X vssd1 vssd1 vccd1 vccd1 _13218_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14195_ _14413_/A vssd1 vssd1 vccd1 vccd1 _14195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10358_ _15515_/Q _10363_/C _10357_/X vssd1 vssd1 vccd1 vccd1 _10360_/C sky130_fd_sc_hd__a21o_1
X_13146_ _14328_/A _13146_/B _13146_/C vssd1 vssd1 vccd1 vccd1 _13149_/B sky130_fd_sc_hd__or3_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _13077_/A _13077_/B _13081_/B vssd1 vssd1 vccd1 vccd1 _15942_/D sky130_fd_sc_hd__nor3_1
X_10289_ _10289_/A vssd1 vssd1 vccd1 vccd1 _10304_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12028_ _15776_/Q _12033_/C _11798_/X vssd1 vssd1 vccd1 vccd1 _12030_/C sky130_fd_sc_hd__a21o_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13979_ _16102_/Q _14117_/B _13979_/C vssd1 vssd1 vccd1 vccd1 _13985_/A sky130_fd_sc_hd__and3_1
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15718_ _15763_/CLK _15718_/D vssd1 vssd1 vccd1 vccd1 _15718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _15655_/CLK _15649_/D vssd1 vssd1 vccd1 vccd1 _15649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ _09168_/Y _09163_/C _09165_/X _09167_/Y vssd1 vssd1 vccd1 vccd1 _09171_/C
+ sky130_fd_sc_hd__a211o_1
X_08121_ _15351_/Q _07734_/B _08120_/Y vssd1 vssd1 vccd1 vccd1 _08242_/B sky130_fd_sc_hd__a21o_2
X_08052_ _08052_/A _08052_/B _08052_/C vssd1 vssd1 vccd1 vccd1 _08053_/B sky130_fd_sc_hd__nand3_1
XFILLER_128_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08954_ _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _08957_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07905_ _16233_/Q _16251_/Q vssd1 vssd1 vccd1 vccd1 _07906_/C sky130_fd_sc_hd__or2_1
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08885_ _08909_/A _08885_/B _08891_/B vssd1 vssd1 vccd1 vccd1 _15285_/D sky130_fd_sc_hd__nor3_1
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07836_ _15863_/Q _15881_/Q vssd1 vssd1 vccd1 vccd1 _08030_/B sky130_fd_sc_hd__xor2_2
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07767_ _12983_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _08083_/A sky130_fd_sc_hd__xnor2_1
XFILLER_112_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09506_ _10663_/A vssd1 vssd1 vccd1 vccd1 _09506_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07698_ _14964_/A _13919_/A _07698_/C vssd1 vssd1 vccd1 vccd1 _07703_/A sky130_fd_sc_hd__and3_1
XFILLER_13_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09437_ _09437_/A vssd1 vssd1 vccd1 vccd1 _15370_/D sky130_fd_sc_hd__clkbuf_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09380_/C vssd1 vssd1 vccd1 vccd1 _09391_/C sky130_fd_sc_hd__clkbuf_1
X_08319_ _08259_/A _08259_/B _08318_/Y vssd1 vssd1 vccd1 vccd1 _08359_/B sky130_fd_sc_hd__a21oi_2
X_09299_ _09306_/B _09299_/B vssd1 vssd1 vccd1 vccd1 _09301_/A sky130_fd_sc_hd__or2_1
X_11330_ _11330_/A vssd1 vssd1 vccd1 vccd1 _15664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11261_ _11268_/B _11261_/B vssd1 vssd1 vccd1 vccd1 _11264_/A sky130_fd_sc_hd__or2_1
X_10212_ input6/X vssd1 vssd1 vccd1 vccd1 _11422_/A sky130_fd_sc_hd__clkbuf_4
X_13000_ _13014_/A _13000_/B _13000_/C vssd1 vssd1 vccd1 vccd1 _13001_/A sky130_fd_sc_hd__and3_1
XFILLER_137_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11192_ _15645_/Q _11198_/C _11137_/X vssd1 vssd1 vccd1 vccd1 _11192_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10143_ _15480_/Q _10199_/B _10143_/C vssd1 vssd1 vccd1 vccd1 _10143_/Y sky130_fd_sc_hd__nand3_1
XFILLER_97_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10074_ _15471_/Q _10074_/B _10074_/C vssd1 vssd1 vccd1 vccd1 _10074_/X sky130_fd_sc_hd__and3_1
X_14951_ _14945_/B _14946_/C _14956_/A _14949_/Y vssd1 vssd1 vccd1 vccd1 _14956_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_121_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13902_ _14402_/A vssd1 vssd1 vccd1 vccd1 _14137_/B sky130_fd_sc_hd__clkbuf_2
X_14882_ _14880_/A _14880_/B _14881_/X vssd1 vssd1 vccd1 vccd1 _16291_/D sky130_fd_sc_hd__a21oi_1
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ _16076_/Q _13832_/C _10950_/C vssd1 vssd1 vccd1 vccd1 _13833_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13764_ _14644_/A _13766_/C vssd1 vssd1 vccd1 vccd1 _13764_/X sky130_fd_sc_hd__or2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10976_ _11204_/A _10979_/C vssd1 vssd1 vccd1 vccd1 _10976_/X sky130_fd_sc_hd__or2_1
XFILLER_71_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15503_ _15512_/CLK _15503_/D vssd1 vssd1 vccd1 vccd1 _15503_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12715_ _15884_/Q _12720_/C _12654_/X vssd1 vssd1 vccd1 vccd1 _12717_/C sky130_fd_sc_hd__a21o_1
X_13695_ _16049_/Q _13794_/B _13701_/C vssd1 vssd1 vccd1 vccd1 _13695_/Y sky130_fd_sc_hd__nand3_1
XFILLER_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15434_ _15483_/CLK _15434_/D vssd1 vssd1 vccd1 vccd1 _15434_/Q sky130_fd_sc_hd__dfxtp_1
X_12646_ _12660_/C vssd1 vssd1 vccd1 vccd1 _12670_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15365_ _15422_/CLK _15365_/D vssd1 vssd1 vccd1 vccd1 _15365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12577_ _12583_/B _12577_/B vssd1 vssd1 vccd1 vccd1 _12579_/A sky130_fd_sc_hd__or2_1
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _14316_/A vssd1 vssd1 vccd1 vccd1 _14316_/X sky130_fd_sc_hd__clkbuf_2
X_11528_ _15696_/Q _11697_/B _11528_/C vssd1 vssd1 vccd1 vccd1 _11528_/Y sky130_fd_sc_hd__nand3_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15296_ _15359_/CLK _15296_/D vssd1 vssd1 vccd1 vccd1 _15296_/Q sky130_fd_sc_hd__dfxtp_1
X_14247_ _16156_/Q _14337_/B _14247_/C vssd1 vssd1 vccd1 vccd1 _14253_/A sky130_fd_sc_hd__and3_1
XFILLER_144_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11459_ _11457_/X _11458_/Y _11454_/B _11455_/C vssd1 vssd1 vccd1 vccd1 _11461_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14178_ _16141_/Q _14185_/C _14177_/X vssd1 vssd1 vccd1 vccd1 _14180_/B sky130_fd_sc_hd__a21oi_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _15952_/Q _13138_/C _14605_/B vssd1 vssd1 vccd1 vccd1 _13129_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08670_ _08670_/A vssd1 vssd1 vccd1 vccd1 _15251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07621_ _13316_/A vssd1 vssd1 vccd1 vccd1 _14901_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ _15337_/Q _09334_/B _09222_/C vssd1 vssd1 vccd1 vccd1 _09222_/Y sky130_fd_sc_hd__nand3_1
XFILLER_10_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09153_ _15328_/Q _09160_/C _08920_/X vssd1 vssd1 vccd1 vccd1 _09153_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08104_ _08104_/A _08224_/A vssd1 vssd1 vccd1 vccd1 _08225_/A sky130_fd_sc_hd__xor2_4
X_09084_ _09096_/C vssd1 vssd1 vccd1 vccd1 _09105_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08035_ _08035_/A _08035_/B vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__xnor2_4
XFILLER_107_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09986_ _10064_/A _09986_/B _09992_/B vssd1 vssd1 vccd1 vccd1 _15455_/D sky130_fd_sc_hd__nor3_1
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08937_ _15294_/Q _09165_/B _08945_/C vssd1 vssd1 vccd1 vccd1 _08937_/X sky130_fd_sc_hd__and3_1
XFILLER_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08868_ _08865_/X _08866_/Y _08867_/Y _08863_/C vssd1 vssd1 vccd1 vccd1 _08870_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07819_ _15872_/Q _07820_/B vssd1 vssd1 vccd1 vccd1 _07821_/A sky130_fd_sc_hd__nand2_1
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08799_ _08799_/A _08799_/B _08799_/C vssd1 vssd1 vccd1 vccd1 _08800_/C sky130_fd_sc_hd__nand3_1
X_10830_ _10830_/A vssd1 vssd1 vccd1 vccd1 _15587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10761_ _15577_/Q _10798_/C _10760_/X vssd1 vssd1 vccd1 vccd1 _10763_/B sky130_fd_sc_hd__a21oi_1
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12500_ _15849_/Q _12554_/B _12500_/C vssd1 vssd1 vccd1 vccd1 _12500_/Y sky130_fd_sc_hd__nand3_1
X_10692_ _10690_/A _10690_/B _10691_/X vssd1 vssd1 vccd1 vccd1 _15564_/D sky130_fd_sc_hd__a21oi_1
X_13480_ _13480_/A _13480_/B _13480_/C vssd1 vssd1 vccd1 vccd1 _13481_/C sky130_fd_sc_hd__nand3_1
XFILLER_13_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12431_ _12431_/A _12431_/B _12431_/C vssd1 vssd1 vccd1 vccd1 _12432_/C sky130_fd_sc_hd__nand3_1
XFILLER_138_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15150_ _15184_/A _15155_/C vssd1 vssd1 vccd1 vccd1 _15150_/Y sky130_fd_sc_hd__nor2_1
X_12362_ _12376_/C vssd1 vssd1 vccd1 vccd1 _12386_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14101_ _14106_/B _14101_/B vssd1 vssd1 vccd1 vccd1 _14103_/A sky130_fd_sc_hd__or2_1
X_11313_ _15662_/Q _11313_/B _11317_/C vssd1 vssd1 vccd1 vccd1 _11313_/Y sky130_fd_sc_hd__nand3_1
X_12293_ _12299_/B _12293_/B vssd1 vssd1 vccd1 vccd1 _12295_/A sky130_fd_sc_hd__or2_1
X_15081_ _15001_/X _15074_/A _15077_/B _15080_/Y vssd1 vssd1 vccd1 vccd1 _16337_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11244_ _15653_/Q _11244_/B _11253_/C vssd1 vssd1 vccd1 vccd1 _11244_/X sky130_fd_sc_hd__and3_1
X_14032_ _16113_/Q _14256_/B _14032_/C vssd1 vssd1 vccd1 vccd1 _14040_/A sky130_fd_sc_hd__and3_1
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11175_ _15643_/Q _11236_/B _11178_/C vssd1 vssd1 vccd1 vccd1 _11175_/X sky130_fd_sc_hd__and3_1
XFILLER_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ _15478_/Q _10239_/B _10135_/C vssd1 vssd1 vccd1 vccd1 _10131_/A sky130_fd_sc_hd__and3_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15983_ _15994_/CLK _15983_/D vssd1 vssd1 vccd1 vccd1 _15983_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10057_ _15475_/Q _15474_/Q _15473_/Q _09831_/X vssd1 vssd1 vccd1 vccd1 _15467_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_57_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14934_ _14814_/X _14932_/A _14933_/Y vssd1 vssd1 vccd1 vccd1 _16304_/D sky130_fd_sc_hd__o21a_1
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14865_ _14866_/B _14866_/C _14866_/A vssd1 vssd1 vccd1 vccd1 _14867_/B sky130_fd_sc_hd__a21o_1
XFILLER_29_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13816_ _13617_/X _13814_/C _13720_/X vssd1 vssd1 vccd1 vccd1 _13816_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_51_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14796_ hold13/A _14795_/C _14718_/X vssd1 vssd1 vccd1 vccd1 _14797_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13747_ _13744_/X _13745_/Y _13746_/Y _13742_/C vssd1 vssd1 vccd1 vccd1 _13749_/B
+ sky130_fd_sc_hd__o211ai_1
X_10959_ _10957_/Y _10953_/C _10955_/X _10956_/Y vssd1 vssd1 vccd1 vccd1 _10960_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ _14073_/A vssd1 vssd1 vccd1 vccd1 _13735_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15417_ _15483_/CLK _15417_/D vssd1 vssd1 vccd1 vccd1 _15417_/Q sky130_fd_sc_hd__dfxtp_1
X_12629_ _12629_/A vssd1 vssd1 vccd1 vccd1 _12861_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15348_ _15348_/CLK _15348_/D vssd1 vssd1 vccd1 vccd1 _15348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15279_ _15359_/CLK _15279_/D vssd1 vssd1 vccd1 vccd1 _15279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _15434_/Q _10010_/B _09847_/C vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__nand3_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09796_/C vssd1 vssd1 vccd1 vccd1 _09811_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _08722_/A vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08653_ _15249_/Q _10965_/C _08657_/C vssd1 vssd1 vccd1 vccd1 _08653_/Y sky130_fd_sc_hd__nand3_1
XFILLER_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07604_ input9/X vssd1 vssd1 vccd1 vccd1 _11898_/A sky130_fd_sc_hd__clkinv_2
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _15240_/Q _10965_/C _08588_/C vssd1 vssd1 vccd1 vccd1 _08584_/Y sky130_fd_sc_hd__nand3_1
XFILLER_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09205_ _09778_/A vssd1 vssd1 vccd1 vccd1 _09205_/X sky130_fd_sc_hd__buf_2
XFILLER_148_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09136_ _09136_/A vssd1 vssd1 vccd1 vccd1 _15323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09067_ _15314_/Q _09067_/B _09067_/C vssd1 vssd1 vccd1 vccd1 _09075_/B sky130_fd_sc_hd__and3_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08018_ _08019_/A _08019_/B vssd1 vssd1 vccd1 vccd1 _08020_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09969_ _09967_/Y _09962_/C _09964_/X _09965_/Y vssd1 vssd1 vccd1 vccd1 _09970_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_58_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12980_ _12980_/A vssd1 vssd1 vccd1 vccd1 _15925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11931_ _15759_/Q _11986_/B _11931_/C vssd1 vssd1 vccd1 vccd1 _11931_/Y sky130_fd_sc_hd__nand3_1
XFILLER_91_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14650_ _14765_/A _14654_/C vssd1 vssd1 vccd1 vccd1 _14652_/A sky130_fd_sc_hd__and2_1
X_11862_ _11862_/A vssd1 vssd1 vccd1 vccd1 _15748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ _16032_/Q _13801_/B _13605_/C vssd1 vssd1 vccd1 vccd1 _13601_/Y sky130_fd_sc_hd__nand3_1
X_10813_ _10825_/C vssd1 vssd1 vccd1 vccd1 _10835_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14581_ _14584_/C vssd1 vssd1 vccd1 vccd1 _14593_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11793_ _15739_/Q _11833_/C _11624_/X vssd1 vssd1 vccd1 vccd1 _11796_/B sky130_fd_sc_hd__a21oi_1
XFILLER_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16320_ _16337_/CLK _16320_/D vssd1 vssd1 vccd1 vccd1 _16320_/Q sky130_fd_sc_hd__dfxtp_1
X_13532_ _13532_/A vssd1 vssd1 vccd1 vccd1 _13738_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10744_ _10744_/A _10744_/B vssd1 vssd1 vccd1 vccd1 _10745_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16251_ _16273_/CLK _16251_/D vssd1 vssd1 vccd1 vccd1 _16251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ _13463_/A vssd1 vssd1 vccd1 vccd1 _16006_/D sky130_fd_sc_hd__clkbuf_1
X_10675_ _10673_/Y _10668_/C _10671_/X _10672_/Y vssd1 vssd1 vccd1 vccd1 _10676_/C
+ sky130_fd_sc_hd__a211o_1
X_15202_ _16359_/CLK _15202_/D vssd1 vssd1 vccd1 vccd1 _15202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12414_ _12583_/A _12414_/B _12414_/C vssd1 vssd1 vccd1 vccd1 _12416_/B sky130_fd_sc_hd__or3_1
X_16182_ _16189_/CLK _16182_/D vssd1 vssd1 vccd1 vccd1 _16182_/Q sky130_fd_sc_hd__dfxtp_2
X_13394_ _15997_/Q _13394_/B _13394_/C vssd1 vssd1 vccd1 vccd1 _13404_/A sky130_fd_sc_hd__and3_1
XFILLER_139_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15133_ _15134_/B _15134_/C _15134_/A vssd1 vssd1 vccd1 vccd1 _15135_/B sky130_fd_sc_hd__a21o_1
X_12345_ _12629_/A vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15064_ _15064_/A _15064_/B _15064_/C vssd1 vssd1 vccd1 vccd1 _15065_/C sky130_fd_sc_hd__nand3_1
XFILLER_142_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12276_ _15815_/Q _12284_/C _12048_/X vssd1 vssd1 vccd1 vccd1 _12276_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14015_ _13925_/X _14011_/B _13926_/X vssd1 vssd1 vccd1 vccd1 _14017_/A sky130_fd_sc_hd__a21oi_1
X_11227_ _11227_/A vssd1 vssd1 vccd1 vccd1 _15649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11158_ _11178_/C vssd1 vssd1 vccd1 vccd1 _11191_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10109_ _10109_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _10111_/B sky130_fd_sc_hd__nor2_1
XFILLER_49_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11089_ _11089_/A _11089_/B vssd1 vssd1 vccd1 vccd1 _11090_/B sky130_fd_sc_hd__nor2_1
X_15966_ _16123_/CLK _15966_/D vssd1 vssd1 vccd1 vccd1 _15966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14917_ _15176_/B vssd1 vssd1 vccd1 vccd1 _14917_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15897_ _07603_/A _15897_/D vssd1 vssd1 vccd1 vccd1 _15897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14848_ _14802_/X _14840_/A _14843_/B _14847_/Y vssd1 vssd1 vccd1 vccd1 _16283_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_24_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14779_ _14825_/A _14779_/B _14785_/A vssd1 vssd1 vccd1 vccd1 _16270_/D sky130_fd_sc_hd__nor3_1
XFILLER_32_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09823_ _10049_/A _09826_/C vssd1 vssd1 vccd1 vccd1 _09823_/X sky130_fd_sc_hd__or2_1
XFILLER_99_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09754_ _15421_/Q _09931_/B _09754_/C vssd1 vssd1 vccd1 vccd1 _09764_/B sky130_fd_sc_hd__and3_1
XFILLER_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08705_ _08705_/A vssd1 vssd1 vccd1 vccd1 _15257_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09685_ _15410_/Q _09740_/B _09692_/C vssd1 vssd1 vccd1 vccd1 _09685_/X sky130_fd_sc_hd__and3_1
XFILLER_66_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk _15584_/CLK vssd1 vssd1 vccd1 vccd1 _15539_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _15247_/Q _08753_/B _08636_/C vssd1 vssd1 vccd1 vccd1 _08636_/Y sky130_fd_sc_hd__nand3_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ hold36/A _08568_/C _12847_/A vssd1 vssd1 vccd1 vccd1 _08567_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08498_ _08498_/A vssd1 vssd1 vccd1 vccd1 _15228_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10460_ _11898_/A vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__buf_4
XFILLER_136_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _15322_/Q _09125_/C _09118_/X vssd1 vssd1 vccd1 vccd1 _09119_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10391_ _15518_/Q _10391_/B _10395_/C vssd1 vssd1 vccd1 vccd1 _10391_/Y sky130_fd_sc_hd__nand3_1
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12130_ _12299_/A _12130_/B _12130_/C vssd1 vssd1 vccd1 vccd1 _12132_/B sky130_fd_sc_hd__or3_1
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12061_ _12629_/A vssd1 vssd1 vccd1 vccd1 _12291_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_89_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11012_ _11012_/A vssd1 vssd1 vccd1 vccd1 _15615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15820_ _07603_/A _15820_/D vssd1 vssd1 vccd1 vccd1 _15820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15751_ _15794_/CLK _15751_/D vssd1 vssd1 vccd1 vccd1 _15751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12963_ _15924_/Q _12968_/C _12855_/X vssd1 vssd1 vccd1 vccd1 _12963_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_84_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15485_/CLK sky130_fd_sc_hd__clkbuf_16
X_14702_ _14901_/A vssd1 vssd1 vccd1 vccd1 _14702_/X sky130_fd_sc_hd__buf_2
X_11914_ _15757_/Q _12025_/B _11923_/C vssd1 vssd1 vccd1 vccd1 _11919_/A sky130_fd_sc_hd__and3_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _15763_/CLK _15682_/D vssd1 vssd1 vccd1 vccd1 _15682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12894_ _15913_/Q _12896_/C _12668_/X vssd1 vssd1 vccd1 vccd1 _12894_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14633_ _14936_/A vssd1 vssd1 vccd1 vccd1 _14716_/A sky130_fd_sc_hd__clkbuf_2
X_11845_ _11883_/A _11845_/B _11845_/C vssd1 vssd1 vccd1 vccd1 _11846_/A sky130_fd_sc_hd__and3_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14562_/A _14562_/B _14561_/Y _14563_/Y vssd1 vssd1 vccd1 vccd1 _16219_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_14_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ _15736_/Q _11774_/C _11775_/X vssd1 vssd1 vccd1 vccd1 _11777_/B sky130_fd_sc_hd__a21oi_1
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16304_/CLK _16303_/D vssd1 vssd1 vccd1 vccd1 _16303_/Q sky130_fd_sc_hd__dfxtp_1
X_13515_ _13515_/A vssd1 vssd1 vccd1 vccd1 _16015_/D sky130_fd_sc_hd__clkbuf_1
X_10727_ _15572_/Q _10895_/B _10734_/C vssd1 vssd1 vccd1 vccd1 _10727_/X sky130_fd_sc_hd__and3_1
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14495_ _14368_/X _14493_/B _14415_/X vssd1 vssd1 vccd1 vccd1 _14495_/Y sky130_fd_sc_hd__a21oi_1
X_16234_ _16247_/CLK _16234_/D vssd1 vssd1 vccd1 vccd1 _16234_/Q sky130_fd_sc_hd__dfxtp_2
X_13446_ _16006_/Q _13451_/C _13342_/X vssd1 vssd1 vccd1 vccd1 _13446_/Y sky130_fd_sc_hd__a21oi_1
X_10658_ _10651_/B _10652_/C _10654_/X _10656_/Y vssd1 vssd1 vccd1 vccd1 _10659_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16165_ _16166_/CLK _16165_/D vssd1 vssd1 vccd1 vccd1 _16165_/Q sky130_fd_sc_hd__dfxtp_1
X_13377_ _13377_/A _13377_/B _13377_/C vssd1 vssd1 vccd1 vccd1 _13378_/C sky130_fd_sc_hd__nand3_1
X_10589_ _10645_/A _10589_/B _10593_/A vssd1 vssd1 vccd1 vccd1 _15549_/D sky130_fd_sc_hd__nor3_1
XFILLER_142_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15116_ _15001_/X _15109_/A _15112_/B _15115_/Y vssd1 vssd1 vccd1 vccd1 _16346_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_127_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12328_ _12326_/Y _12321_/C _12323_/X _12324_/Y vssd1 vssd1 vccd1 vccd1 _12329_/C
+ sky130_fd_sc_hd__a211o_1
X_16096_ _16103_/CLK _16096_/D vssd1 vssd1 vccd1 vccd1 _16096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15047_ _15152_/A _15051_/C vssd1 vssd1 vccd1 vccd1 _15049_/A sky130_fd_sc_hd__and2_1
X_12259_ _12259_/A _12259_/B _12259_/C vssd1 vssd1 vccd1 vccd1 _12260_/C sky130_fd_sc_hd__nand3_1
XFILLER_68_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15949_ _16100_/CLK _15949_/D vssd1 vssd1 vccd1 vccd1 _15949_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_75_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15339_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09470_ _09470_/A _09470_/B vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__nor2_1
X_08421_ _08421_/A _08421_/B _08421_/C vssd1 vssd1 vccd1 vccd1 _15215_/D sky130_fd_sc_hd__nor3_4
XFILLER_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08352_ _08352_/A _08304_/A vssd1 vssd1 vccd1 vccd1 _08356_/B sky130_fd_sc_hd__or2b_1
XFILLER_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08283_ _08283_/A _08267_/A vssd1 vssd1 vccd1 vccd1 _08283_/X sky130_fd_sc_hd__or2b_1
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09806_ _09804_/Y _09799_/C _09802_/X _09803_/Y vssd1 vssd1 vccd1 vccd1 _09807_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07998_ _07999_/A _07999_/B vssd1 vssd1 vccd1 vccd1 _08209_/A sky130_fd_sc_hd__nand2_2
X_09737_ _09735_/Y _09731_/C _09733_/X _09734_/Y vssd1 vssd1 vccd1 vccd1 _09738_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_66_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15274_/CLK sky130_fd_sc_hd__clkbuf_16
X_09668_ _09668_/A _09668_/B _09668_/C vssd1 vssd1 vccd1 vccd1 _09669_/C sky130_fd_sc_hd__nand3_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _08619_/A _08619_/B _08619_/C vssd1 vssd1 vccd1 vccd1 _08620_/C sky130_fd_sc_hd__nand3_1
XFILLER_131_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09599_ _09599_/A vssd1 vssd1 vccd1 vccd1 _15394_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11631_/B _11631_/C _11631_/A vssd1 vssd1 vccd1 vccd1 _11632_/B sky130_fd_sc_hd__a21o_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11561_ _15709_/Q _15708_/Q _15707_/Q _11560_/X vssd1 vssd1 vccd1 vccd1 _15701_/D
+ sky130_fd_sc_hd__o31a_1
X_13300_ _13300_/A _13300_/B vssd1 vssd1 vccd1 vccd1 _13301_/B sky130_fd_sc_hd__nor2_1
X_10512_ _15538_/Q _10512_/B _10512_/C vssd1 vssd1 vccd1 vccd1 _10520_/B sky130_fd_sc_hd__and3_1
XFILLER_109_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14280_ _14195_/X _14277_/B _14279_/Y vssd1 vssd1 vccd1 vccd1 _16159_/D sky130_fd_sc_hd__o21a_1
X_11492_ _11492_/A _11492_/B vssd1 vssd1 vccd1 vccd1 _11497_/C sky130_fd_sc_hd__nor2_1
XFILLER_7_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13231_ _13231_/A vssd1 vssd1 vccd1 vccd1 _15966_/D sky130_fd_sc_hd__clkbuf_1
X_10443_ _10441_/Y _10437_/C _10439_/X _10440_/Y vssd1 vssd1 vccd1 vccd1 _10444_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13162_ _15957_/Q _14379_/A _13162_/C vssd1 vssd1 vccd1 vccd1 _13169_/A sky130_fd_sc_hd__and3_1
XFILLER_108_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10374_ _15517_/Q _10375_/C _10373_/X vssd1 vssd1 vccd1 vccd1 _10374_/Y sky130_fd_sc_hd__a21oi_1
X_12113_ _12113_/A vssd1 vssd1 vccd1 vccd1 _15787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13093_ _13109_/C vssd1 vssd1 vccd1 vccd1 _13127_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12044_ _12042_/Y _12037_/C _12039_/X _12040_/Y vssd1 vssd1 vccd1 vccd1 _12045_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15803_ _07603_/A _15803_/D vssd1 vssd1 vccd1 vccd1 _15803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13995_ _14261_/A vssd1 vssd1 vccd1 vccd1 _14221_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _16327_/CLK sky130_fd_sc_hd__clkbuf_16
X_15734_ _15763_/CLK _15734_/D vssd1 vssd1 vccd1 vccd1 _15734_/Q sky130_fd_sc_hd__dfxtp_1
X_12946_ _12946_/A vssd1 vssd1 vccd1 vccd1 _15920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15665_ _15665_/CLK _15665_/D vssd1 vssd1 vccd1 vccd1 _15665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12877_ _12908_/C vssd1 vssd1 vccd1 vccd1 _12914_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _13921_/X _14612_/B _14615_/Y vssd1 vssd1 vccd1 vccd1 _16231_/D sky130_fd_sc_hd__o21a_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _15744_/Q _11833_/C _11713_/X vssd1 vssd1 vccd1 vccd1 _11828_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15596_ _15194_/Q _15596_/D vssd1 vssd1 vccd1 vccd1 _15596_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14626_/A _14547_/B _14551_/A vssd1 vssd1 vccd1 vccd1 _16216_/D sky130_fd_sc_hd__nor3_1
X_11759_ _15734_/Q _11819_/B _11767_/C vssd1 vssd1 vccd1 vccd1 _11759_/X sky130_fd_sc_hd__and3_1
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14478_ _14517_/A _14478_/B _14481_/B vssd1 vssd1 vccd1 vccd1 _16200_/D sky130_fd_sc_hd__nor3_1
X_16217_ _16240_/CLK _16217_/D vssd1 vssd1 vccd1 vccd1 _16217_/Q sky130_fd_sc_hd__dfxtp_2
X_13429_ _13429_/A vssd1 vssd1 vccd1 vccd1 _16001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16148_ _16148_/CLK _16148_/D vssd1 vssd1 vccd1 vccd1 _16148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08970_ _15299_/Q _09008_/C _08735_/X vssd1 vssd1 vccd1 vccd1 _08972_/B sky130_fd_sc_hd__a21oi_1
X_16079_ _16124_/CLK _16079_/D vssd1 vssd1 vccd1 vccd1 _16079_/Q sky130_fd_sc_hd__dfxtp_1
X_07921_ _15602_/Q _07954_/B vssd1 vssd1 vccd1 vccd1 _07922_/B sky130_fd_sc_hd__xnor2_2
XFILLER_102_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07852_ _16044_/Q vssd1 vssd1 vccd1 vccd1 _13729_/C sky130_fd_sc_hd__clkinv_4
Xinput1 in1[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07783_ _15710_/Q _07783_/B vssd1 vssd1 vccd1 vccd1 _07784_/B sky130_fd_sc_hd__or2_1
XFILLER_110_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16264_/CLK sky130_fd_sc_hd__clkbuf_16
X_09522_ _15384_/Q _09577_/B _09522_/C vssd1 vssd1 vccd1 vccd1 _09531_/A sky130_fd_sc_hd__and3_1
XFILLER_83_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09453_ _10610_/A vssd1 vssd1 vccd1 vccd1 _09453_/X sky130_fd_sc_hd__buf_2
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08404_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08404_/X sky130_fd_sc_hd__and2_1
X_09384_ _09401_/A _09384_/B _09384_/C vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__and3_1
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08335_ _15086_/A vssd1 vssd1 vccd1 vccd1 _08335_/X sky130_fd_sc_hd__clkbuf_4
X_08266_ _08266_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08283_/A sky130_fd_sc_hd__xnor2_2
X_08197_ _08287_/A _08287_/B vssd1 vssd1 vccd1 vccd1 _08198_/B sky130_fd_sc_hd__xor2_2
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10090_ input5/X vssd1 vssd1 vccd1 vccd1 _11303_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_39_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16142_/CLK sky130_fd_sc_hd__clkbuf_16
X_12800_ _13847_/A vssd1 vssd1 vccd1 vccd1 _13018_/B sky130_fd_sc_hd__buf_2
X_13780_ _16066_/Q _13785_/C _07634_/A vssd1 vssd1 vccd1 vccd1 _13782_/C sky130_fd_sc_hd__a21o_1
XFILLER_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10992_ _11569_/A vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _12729_/Y _12724_/C _12727_/X _12728_/Y vssd1 vssd1 vccd1 vccd1 _12732_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _15483_/CLK _15450_/D vssd1 vssd1 vccd1 vccd1 _15450_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _15876_/Q _12670_/C _12661_/X vssd1 vssd1 vccd1 vccd1 _12662_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14398_/B _14397_/Y _14398_/A vssd1 vssd1 vccd1 vccd1 _14401_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11842_/A vssd1 vssd1 vccd1 vccd1 _11653_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15484_/CLK _15381_/D vssd1 vssd1 vccd1 vccd1 _15381_/Q sky130_fd_sc_hd__dfxtp_1
X_12593_ _15865_/Q _12593_/B _12601_/C vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__and3_1
XFILLER_129_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14332_ _14434_/A vssd1 vssd1 vccd1 vccd1 _14427_/A sky130_fd_sc_hd__clkbuf_2
X_11544_ _11550_/A _11542_/Y _11543_/Y _11538_/C vssd1 vssd1 vccd1 vccd1 _11546_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _16159_/Q _14269_/C _14177_/X vssd1 vssd1 vccd1 vccd1 _14265_/B sky130_fd_sc_hd__a21oi_1
X_11475_ _11471_/X _11473_/Y _11474_/Y _11469_/C vssd1 vssd1 vccd1 vccd1 _11477_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_143_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371__20 vssd1 vssd1 vccd1 vccd1 _16371__20/HI io_oeb[3] sky130_fd_sc_hd__conb_1
X_16002_ _16011_/CLK _16002_/D vssd1 vssd1 vccd1 vccd1 _16002_/Q sky130_fd_sc_hd__dfxtp_1
X_13214_ _13240_/C vssd1 vssd1 vccd1 vccd1 _13246_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10426_ _15525_/Q _10654_/B _10426_/C vssd1 vssd1 vccd1 vccd1 _10426_/X sky130_fd_sc_hd__and3_1
XFILLER_124_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14194_ _14190_/X _14192_/B _14193_/Y vssd1 vssd1 vccd1 vccd1 _16140_/D sky130_fd_sc_hd__o21a_1
X_13145_ _13715_/A vssd1 vssd1 vccd1 vccd1 _14328_/A sky130_fd_sc_hd__buf_2
X_10357_ _11222_/A vssd1 vssd1 vccd1 vccd1 _10357_/X sky130_fd_sc_hd__clkbuf_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _13074_/Y _13069_/C _13081_/A _13072_/Y vssd1 vssd1 vccd1 vccd1 _13081_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_112_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10288_ _15511_/Q _15510_/Q _15509_/Q _10119_/X vssd1 vssd1 vccd1 vccd1 _15503_/D
+ sky130_fd_sc_hd__o31a_1
X_12027_ _15776_/Q _12085_/B _12033_/C vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__nand3_1
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13978_ _16102_/Q _14003_/C _13822_/X vssd1 vssd1 vccd1 vccd1 _13980_/B sky130_fd_sc_hd__a21oi_1
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15717_ _15763_/CLK _15717_/D vssd1 vssd1 vccd1 vccd1 _15717_/Q sky130_fd_sc_hd__dfxtp_1
X_12929_ _12941_/C vssd1 vssd1 vccd1 vccd1 _12949_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15648_ _15655_/CLK _15648_/D vssd1 vssd1 vccd1 vccd1 _15648_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15579_ _15194_/Q _15579_/D vssd1 vssd1 vccd1 vccd1 _15579_/Q sky130_fd_sc_hd__dfxtp_1
X_08120_ _09256_/A _09138_/A vssd1 vssd1 vccd1 vccd1 _08120_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08051_ _08052_/A _08052_/B _08052_/C vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__a21o_1
XFILLER_119_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08953_ _08961_/B _08953_/B vssd1 vssd1 vccd1 vccd1 _08957_/A sky130_fd_sc_hd__or2_1
XFILLER_130_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07904_ _16233_/Q _16251_/Q vssd1 vssd1 vccd1 vccd1 _07963_/A sky130_fd_sc_hd__nand2_2
XFILLER_57_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08884_ _08882_/Y _08878_/C _08891_/A _08881_/Y vssd1 vssd1 vccd1 vccd1 _08891_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07835_ _16134_/Q vssd1 vssd1 vccd1 vccd1 _14207_/C sky130_fd_sc_hd__clkinv_4
XFILLER_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07766_ _08098_/A _07766_/B vssd1 vssd1 vccd1 vccd1 _07767_/B sky130_fd_sc_hd__xnor2_4
XFILLER_65_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09505_ _10947_/A vssd1 vssd1 vccd1 vccd1 _10663_/A sky130_fd_sc_hd__buf_4
XFILLER_65_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07697_ _15050_/A vssd1 vssd1 vccd1 vccd1 _13919_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ _09458_/A _09436_/B _09436_/C vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__and3_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09367_/A vssd1 vssd1 vccd1 vccd1 _09380_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_21_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08318_ _08318_/A _08318_/B vssd1 vssd1 vccd1 vccd1 _08318_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09298_ _15350_/Q _09297_/C _09180_/X vssd1 vssd1 vccd1 vccd1 _09299_/B sky130_fd_sc_hd__a21oi_1
X_08249_ _08249_/A _08249_/B _08249_/C vssd1 vssd1 vccd1 vccd1 _08250_/B sky130_fd_sc_hd__and3_1
XFILLER_119_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ _15655_/Q _11259_/C _11199_/X vssd1 vssd1 vccd1 vccd1 _11261_/B sky130_fd_sc_hd__a21oi_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10211_ _10211_/A vssd1 vssd1 vccd1 vccd1 _15490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11191_ _15645_/Q _11367_/B _11191_/C vssd1 vssd1 vccd1 vccd1 _11202_/A sky130_fd_sc_hd__and3_1
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10142_ _15481_/Q _10143_/C _10083_/X vssd1 vssd1 vccd1 vccd1 _10142_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ _10073_/A vssd1 vssd1 vccd1 vccd1 _15469_/D sky130_fd_sc_hd__clkbuf_1
X_14950_ _14956_/A _14949_/Y _14945_/B _14946_/C vssd1 vssd1 vccd1 vccd1 _14952_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13901_ _13896_/B _13895_/Y _13896_/A vssd1 vssd1 vccd1 vccd1 _13901_/Y sky130_fd_sc_hd__o21bai_1
X_14881_ _15041_/A _14881_/B vssd1 vssd1 vccd1 vccd1 _14881_/X sky130_fd_sc_hd__or2_1
X_13832_ _16076_/Q _14080_/B _13832_/C vssd1 vssd1 vccd1 vccd1 _13832_/X sky130_fd_sc_hd__and3_1
XFILLER_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13763_ _13763_/A _13763_/B vssd1 vssd1 vccd1 vccd1 _13766_/C sky130_fd_sc_hd__nor2_1
XFILLER_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10975_ _10975_/A _10975_/B vssd1 vssd1 vccd1 vccd1 _10979_/C sky130_fd_sc_hd__nor2_1
XFILLER_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _15224_/Q _15502_/D vssd1 vssd1 vccd1 vccd1 _15502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12714_ _15884_/Q _12935_/B _12720_/C vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__nand3_1
XFILLER_31_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13694_ _16050_/Q _13701_/C _13693_/X vssd1 vssd1 vccd1 vccd1 _13694_/Y sky130_fd_sc_hd__a21oi_1
X_15433_ _15483_/CLK _15433_/D vssd1 vssd1 vccd1 vccd1 _15433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12645_ _15872_/Q vssd1 vssd1 vccd1 vccd1 _12660_/C sky130_fd_sc_hd__inv_2
XFILLER_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15364_ _15377_/CLK _15364_/D vssd1 vssd1 vccd1 vccd1 _15364_/Q sky130_fd_sc_hd__dfxtp_1
X_12576_ _15862_/Q _12575_/C _12347_/X vssd1 vssd1 vccd1 vccd1 _12577_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14315_ _14313_/X _14315_/B vssd1 vssd1 vccd1 vccd1 _14315_/X sky130_fd_sc_hd__and2b_1
X_11527_ _15697_/Q _11528_/C _11526_/X vssd1 vssd1 vccd1 vccd1 _11527_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_144_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15295_ _15359_/CLK _15295_/D vssd1 vssd1 vccd1 vccd1 _15295_/Q sky130_fd_sc_hd__dfxtp_1
X_14246_ _16156_/Q _14269_/C _14069_/X vssd1 vssd1 vccd1 vccd1 _14248_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11458_ _15687_/Q _11466_/C _11230_/X vssd1 vssd1 vccd1 vccd1 _11458_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10409_ _10983_/A vssd1 vssd1 vccd1 vccd1 _10409_/X sky130_fd_sc_hd__clkbuf_2
X_14177_ _14395_/A vssd1 vssd1 vccd1 vccd1 _14177_/X sky130_fd_sc_hd__clkbuf_2
X_11389_ _11401_/C vssd1 vssd1 vccd1 vccd1 _11409_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13847_/A vssd1 vssd1 vccd1 vccd1 _14605_/B sky130_fd_sc_hd__clkbuf_4
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _15940_/Q _14031_/A _13059_/C vssd1 vssd1 vccd1 vccd1 _13059_/Y sky130_fd_sc_hd__nand3_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ _15021_/A vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09221_ _15338_/Q _09222_/C _09220_/X vssd1 vssd1 vccd1 vccd1 _09221_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _15328_/Q _09211_/B _09152_/C vssd1 vssd1 vccd1 vccd1 _09152_/X sky130_fd_sc_hd__and3_1
XFILLER_147_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08103_ _08103_/A _08103_/B vssd1 vssd1 vccd1 vccd1 _08224_/A sky130_fd_sc_hd__xnor2_4
X_09083_ _15306_/Q vssd1 vssd1 vccd1 vccd1 _09096_/C sky130_fd_sc_hd__inv_2
X_08034_ _08034_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08035_/B sky130_fd_sc_hd__nor2_2
XFILLER_116_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09985_ _09983_/Y _09977_/C _09992_/A _09982_/Y vssd1 vssd1 vccd1 vccd1 _09992_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_89_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08936_ _09801_/A vssd1 vssd1 vccd1 vccd1 _09165_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08867_ _15283_/Q _09047_/B _08867_/C vssd1 vssd1 vccd1 vccd1 _08867_/Y sky130_fd_sc_hd__nand3_1
XFILLER_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07818_ _07818_/A _07818_/B vssd1 vssd1 vccd1 vccd1 _07820_/B sky130_fd_sc_hd__xor2_1
X_08798_ _08799_/B _08799_/C _08799_/A vssd1 vssd1 vccd1 vccd1 _08800_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07749_ _15449_/Q _15431_/Q vssd1 vssd1 vccd1 vccd1 _07750_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10760_ _11624_/A vssd1 vssd1 vccd1 vccd1 _10760_/X sky130_fd_sc_hd__buf_2
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09419_ _09419_/A _09419_/B _09419_/C vssd1 vssd1 vccd1 vccd1 _09421_/B sky130_fd_sc_hd__or3_1
X_10691_ _10916_/A _10694_/C vssd1 vssd1 vccd1 vccd1 _10691_/X sky130_fd_sc_hd__or2_1
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12430_ _12431_/B _12431_/C _12431_/A vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__a21o_1
XFILLER_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12361_ _12361_/A vssd1 vssd1 vccd1 vccd1 _12376_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14100_ _16124_/Q _14099_/C _13708_/X vssd1 vssd1 vccd1 vccd1 _14101_/B sky130_fd_sc_hd__a21oi_1
X_11312_ _15663_/Q _11317_/C _11137_/X vssd1 vssd1 vccd1 vccd1 _11312_/Y sky130_fd_sc_hd__a21oi_1
X_15080_ _15184_/A _15085_/C vssd1 vssd1 vccd1 vccd1 _15080_/Y sky130_fd_sc_hd__nor2_1
X_12292_ _15817_/Q _12291_/C _12063_/X vssd1 vssd1 vccd1 vccd1 _12293_/B sky130_fd_sc_hd__a21oi_1
X_14031_ _14031_/A vssd1 vssd1 vccd1 vccd1 _14256_/B sky130_fd_sc_hd__buf_2
X_11243_ _11243_/A vssd1 vssd1 vccd1 vccd1 _15651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11174_ _11174_/A vssd1 vssd1 vccd1 vccd1 _15641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ _15478_/Q _10162_/C _09893_/X vssd1 vssd1 vccd1 vccd1 _10127_/B sky130_fd_sc_hd__a21oi_1
X_15982_ _15984_/CLK _15982_/D vssd1 vssd1 vccd1 vccd1 _15982_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10056_ _10056_/A vssd1 vssd1 vccd1 vccd1 _15466_/D sky130_fd_sc_hd__clkbuf_1
X_14933_ _14772_/X _14932_/A _14815_/X vssd1 vssd1 vccd1 vccd1 _14933_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14864_ _16293_/Q _14863_/C _14744_/X vssd1 vssd1 vccd1 vccd1 _14866_/C sky130_fd_sc_hd__a21o_1
XFILLER_29_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13815_ _13815_/A vssd1 vssd1 vccd1 vccd1 _16069_/D sky130_fd_sc_hd__clkbuf_1
X_14795_ hold13/A _14953_/B _14795_/C vssd1 vssd1 vccd1 vccd1 _14797_/A sky130_fd_sc_hd__and3_1
X_13746_ _16058_/Q _13794_/B _13752_/C vssd1 vssd1 vccd1 vccd1 _13746_/Y sky130_fd_sc_hd__nand3_1
XFILLER_44_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10958_ _10955_/X _10956_/Y _10957_/Y _10953_/C vssd1 vssd1 vccd1 vccd1 _10960_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_71_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13677_ _14163_/A vssd1 vssd1 vccd1 vccd1 _14073_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10889_ _15598_/Q _10890_/C _10663_/X vssd1 vssd1 vccd1 vccd1 _10889_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_148_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15416_ _15483_/CLK _15416_/D vssd1 vssd1 vccd1 vccd1 _15416_/Q sky130_fd_sc_hd__dfxtp_1
X_12628_ _12652_/A _12628_/B _12634_/B vssd1 vssd1 vccd1 vccd1 _15869_/D sky130_fd_sc_hd__nor3_1
XFILLER_8_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15347_ _15348_/CLK _15347_/D vssd1 vssd1 vccd1 vccd1 _15347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ _15860_/Q _12675_/B _12568_/C vssd1 vssd1 vccd1 vccd1 _12559_/X sky130_fd_sc_hd__and3_1
XFILLER_129_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15278_ _15359_/CLK _15278_/D vssd1 vssd1 vccd1 vccd1 _15278_/Q sky130_fd_sc_hd__dfxtp_1
X_14229_ _16151_/Q _14228_/C _14004_/X vssd1 vssd1 vccd1 vccd1 _14230_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09784_/C vssd1 vssd1 vccd1 vccd1 _09796_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08721_ _08719_/A _08719_/B _08720_/X vssd1 vssd1 vccd1 vccd1 _15259_/D sky130_fd_sc_hd__a21oi_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08652_ _15250_/Q _08657_/C _08524_/X vssd1 vssd1 vccd1 vccd1 _08652_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07603_ _07603_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _15196_/D sky130_fd_sc_hd__nor2_1
X_08583_ _15241_/Q _08588_/C _08524_/X vssd1 vssd1 vccd1 vccd1 _08583_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09204_ _15336_/Q _09432_/B _09211_/C vssd1 vssd1 vccd1 vccd1 _09208_/B sky130_fd_sc_hd__nand3_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09135_ _09171_/A _09135_/B _09135_/C vssd1 vssd1 vccd1 vccd1 _09136_/A sky130_fd_sc_hd__and3_1
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09066_ _09066_/A _09066_/B _09070_/B vssd1 vssd1 vccd1 vccd1 _15312_/D sky130_fd_sc_hd__nor3_1
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08017_ _12304_/A _07869_/B _08016_/X vssd1 vssd1 vccd1 vccd1 _08019_/B sky130_fd_sc_hd__o21a_1
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09968_ _09964_/X _09965_/Y _09967_/Y _09962_/C vssd1 vssd1 vccd1 vccd1 _09970_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08919_ _15292_/Q _08919_/B _08919_/C vssd1 vssd1 vccd1 vccd1 _08919_/X sky130_fd_sc_hd__and3_1
XFILLER_58_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09899_ _09900_/B _09900_/C _09900_/A vssd1 vssd1 vccd1 vccd1 _09901_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11930_ _15760_/Q _11931_/C _11812_/X vssd1 vssd1 vccd1 vccd1 _11930_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11861_ _11883_/A _11861_/B _11861_/C vssd1 vssd1 vccd1 vccd1 _11862_/A sky130_fd_sc_hd__and3_1
XFILLER_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13600_ _14395_/A vssd1 vssd1 vccd1 vccd1 _13801_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10812_ _10812_/A vssd1 vssd1 vccd1 vccd1 _10825_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14580_ hold26/X hold23/X hold27/X _14421_/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__o31a_2
X_11792_ _11827_/C vssd1 vssd1 vccd1 vccd1 _11833_/C sky130_fd_sc_hd__clkbuf_2
X_13531_ _13531_/A vssd1 vssd1 vccd1 vccd1 _16019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10743_ _10750_/B _10743_/B vssd1 vssd1 vccd1 vccd1 _10745_/A sky130_fd_sc_hd__or2_1
XFILLER_43_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16250_ _16268_/CLK _16250_/D vssd1 vssd1 vccd1 vccd1 _16250_/Q sky130_fd_sc_hd__dfxtp_1
X_13462_ _13481_/A _13462_/B _13462_/C vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__and3_1
X_10674_ _10671_/X _10672_/Y _10673_/Y _10668_/C vssd1 vssd1 vccd1 vccd1 _10676_/B
+ sky130_fd_sc_hd__o211ai_1
X_15201_ _16241_/CLK _15201_/D vssd1 vssd1 vccd1 vccd1 _15201_/Q sky130_fd_sc_hd__dfxtp_2
X_12413_ _12413_/A vssd1 vssd1 vccd1 vccd1 _12454_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16181_ _16189_/CLK _16181_/D vssd1 vssd1 vccd1 vccd1 _16181_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13393_ _13393_/A vssd1 vssd1 vccd1 vccd1 _15994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15132_ _16356_/Q _15131_/C _13981_/B vssd1 vssd1 vccd1 vccd1 _15134_/C sky130_fd_sc_hd__a21o_1
X_12344_ _12368_/A _12344_/B _12350_/B vssd1 vssd1 vccd1 vccd1 _15824_/D sky130_fd_sc_hd__nor3_1
XFILLER_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15063_ _15064_/B _15064_/C _15064_/A vssd1 vssd1 vccd1 vccd1 _15065_/B sky130_fd_sc_hd__a21o_1
XFILLER_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12275_ _15815_/Q _12391_/B _12284_/C vssd1 vssd1 vccd1 vccd1 _12275_/X sky130_fd_sc_hd__and3_1
XFILLER_141_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14014_ _13920_/X _14011_/B _14013_/Y vssd1 vssd1 vccd1 vccd1 _16105_/D sky130_fd_sc_hd__o21a_1
X_11226_ _11249_/A _11226_/B _11226_/C vssd1 vssd1 vccd1 vccd1 _11227_/A sky130_fd_sc_hd__and3_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11157_ _11169_/C vssd1 vssd1 vccd1 vccd1 _11178_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10108_ _10115_/B _10108_/B vssd1 vssd1 vccd1 vccd1 _10111_/A sky130_fd_sc_hd__or2_1
XFILLER_67_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11088_ _11094_/B _11088_/B vssd1 vssd1 vccd1 vccd1 _11090_/A sky130_fd_sc_hd__or2_1
X_15965_ _16119_/CLK _15965_/D vssd1 vssd1 vccd1 vccd1 _15965_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10039_ _15464_/Q _10102_/B _10043_/C vssd1 vssd1 vccd1 vccd1 _10039_/Y sky130_fd_sc_hd__nand3_1
XFILLER_82_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14916_ hold17/X _14953_/B _14916_/C vssd1 vssd1 vccd1 vccd1 _14919_/A sky130_fd_sc_hd__and3_1
XFILLER_64_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15896_ _07603_/A _15896_/D vssd1 vssd1 vccd1 vccd1 _15896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14847_ _14847_/A _14853_/C vssd1 vssd1 vccd1 vccd1 _14847_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14778_ _16274_/Q _14778_/B _14782_/C vssd1 vssd1 vccd1 vccd1 _14785_/A sky130_fd_sc_hd__and3_1
XFILLER_32_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13729_ _16056_/Q _14071_/B _13729_/C vssd1 vssd1 vccd1 vccd1 _13734_/A sky130_fd_sc_hd__and3_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09822_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09826_/C sky130_fd_sc_hd__nor2_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09753_ _09775_/A _09753_/B _09758_/B vssd1 vssd1 vccd1 vccd1 _15419_/D sky130_fd_sc_hd__nor3_1
X_08704_ _08704_/A _08704_/B _08704_/C vssd1 vssd1 vccd1 vccd1 _08705_/A sky130_fd_sc_hd__and3_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09684_ _09684_/A vssd1 vssd1 vccd1 vccd1 _15408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08635_ _15248_/Q _08636_/C _08634_/X vssd1 vssd1 vccd1 vccd1 _08635_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ hold36/A _11128_/A _08568_/C vssd1 vssd1 vccd1 vccd1 _08566_/X sky130_fd_sc_hd__and3_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08497_ _08519_/A _08497_/B _08497_/C vssd1 vssd1 vccd1 vccd1 _08498_/A sky130_fd_sc_hd__and3_1
XFILLER_120_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09118_ _09693_/A vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__buf_2
X_10390_ _15519_/Q _10395_/C _10269_/X vssd1 vssd1 vccd1 vccd1 _10390_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09049_ _09047_/Y _09043_/C _09045_/X _09046_/Y vssd1 vssd1 vccd1 vccd1 _09050_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _12084_/A _12060_/B _12066_/B vssd1 vssd1 vccd1 vccd1 _15779_/D sky130_fd_sc_hd__nor3_1
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11011_ _11019_/A _11011_/B _11011_/C vssd1 vssd1 vccd1 vccd1 _11012_/A sky130_fd_sc_hd__and3_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15750_ _15794_/CLK _15750_/D vssd1 vssd1 vccd1 vccd1 _15750_/Q sky130_fd_sc_hd__dfxtp_1
X_12962_ _15924_/Q _13071_/B _12962_/C vssd1 vssd1 vccd1 vccd1 _12971_/A sky130_fd_sc_hd__and3_1
XFILLER_46_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11913_ _15757_/Q _11950_/C _11912_/X vssd1 vssd1 vccd1 vccd1 _11915_/B sky130_fd_sc_hd__a21oi_1
X_14701_ _14706_/C vssd1 vssd1 vccd1 vccd1 _14717_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _15763_/CLK _15681_/D vssd1 vssd1 vccd1 vccd1 _15681_/Q sky130_fd_sc_hd__dfxtp_1
X_12893_ _15913_/Q _12947_/B _12896_/C vssd1 vssd1 vccd1 vccd1 _12893_/X sky130_fd_sc_hd__and3_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11844_ _11843_/B _11843_/C _11615_/X vssd1 vssd1 vccd1 vccd1 _11845_/C sky130_fd_sc_hd__o21ai_1
X_14632_ _14632_/A vssd1 vssd1 vccd1 vccd1 _16235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14562_/X _14561_/Y _14648_/A vssd1 vssd1 vccd1 vccd1 _14563_/Y sky130_fd_sc_hd__a21oi_1
X_11775_ _12631_/A vssd1 vssd1 vccd1 vccd1 _11775_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16304_/CLK _16302_/D vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _10726_/A vssd1 vssd1 vccd1 vccd1 _15570_/D sky130_fd_sc_hd__clkbuf_1
X_13514_ _13538_/A _13514_/B _13514_/C vssd1 vssd1 vccd1 vccd1 _13515_/A sky130_fd_sc_hd__and3_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14494_ _14408_/X _14492_/B _14493_/Y vssd1 vssd1 vccd1 vccd1 _16203_/D sky130_fd_sc_hd__o21a_1
X_16233_ _16268_/CLK _16233_/D vssd1 vssd1 vccd1 vccd1 _16233_/Q sky130_fd_sc_hd__dfxtp_1
X_13445_ _16006_/Q _13648_/B _13445_/C vssd1 vssd1 vccd1 vccd1 _13455_/A sky130_fd_sc_hd__and3_1
X_10657_ _10654_/X _10656_/Y _10651_/B _10652_/C vssd1 vssd1 vccd1 vccd1 _10659_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16164_ _16187_/CLK _16164_/D vssd1 vssd1 vccd1 vccd1 _16164_/Q sky130_fd_sc_hd__dfxtp_2
X_13376_ _13377_/B _13377_/C _13377_/A vssd1 vssd1 vccd1 vccd1 _13378_/B sky130_fd_sc_hd__a21o_1
X_10588_ _15550_/Q _10817_/B _10596_/C vssd1 vssd1 vccd1 vccd1 _10593_/A sky130_fd_sc_hd__and3_1
XFILLER_127_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15115_ _15184_/A _15120_/C vssd1 vssd1 vccd1 vccd1 _15115_/Y sky130_fd_sc_hd__nor2_1
X_12327_ _12323_/X _12324_/Y _12326_/Y _12321_/C vssd1 vssd1 vccd1 vccd1 _12329_/B
+ sky130_fd_sc_hd__o211ai_1
X_16095_ _16103_/CLK _16095_/D vssd1 vssd1 vccd1 vccd1 _16095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15046_ _15001_/X _15038_/A _15041_/B _15045_/Y vssd1 vssd1 vccd1 vccd1 _16328_/D
+ sky130_fd_sc_hd__o31a_1
X_12258_ _12259_/B _12259_/C _12259_/A vssd1 vssd1 vccd1 vccd1 _12260_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11209_ _11208_/B _11208_/C _11038_/X vssd1 vssd1 vccd1 vccd1 _11210_/C sky130_fd_sc_hd__o21ai_1
XFILLER_96_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ _12187_/B _12187_/C _12188_/X vssd1 vssd1 vccd1 vccd1 _12190_/C sky130_fd_sc_hd__o21ai_1
XFILLER_96_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15948_ _15956_/CLK _15948_/D vssd1 vssd1 vccd1 vccd1 _15948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15879_ _15907_/CLK _15879_/D vssd1 vssd1 vccd1 vccd1 _15879_/Q sky130_fd_sc_hd__dfxtp_1
X_08420_ _08420_/A spike_out[0] _08420_/C vssd1 vssd1 vccd1 vccd1 _08421_/C sky130_fd_sc_hd__nor3_2
XFILLER_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08356_/A sky130_fd_sc_hd__or2_1
XFILLER_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08282_ _08282_/A _08268_/A vssd1 vssd1 vccd1 vccd1 _08365_/A sky130_fd_sc_hd__or2b_2
XFILLER_149_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09805_ _09802_/X _09803_/Y _09804_/Y _09799_/C vssd1 vssd1 vccd1 vccd1 _09807_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_87_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07997_ _14161_/C _14247_/C _07996_/Y vssd1 vssd1 vccd1 vccd1 _07999_/B sky130_fd_sc_hd__o21ai_2
XFILLER_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09736_ _09733_/X _09734_/Y _09735_/Y _09731_/C vssd1 vssd1 vccd1 vccd1 _09738_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ _09668_/B _09668_/C _09668_/A vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _08619_/B _08619_/C _08619_/A vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09635_/A _09598_/B _09598_/C vssd1 vssd1 vccd1 vccd1 _09599_/A sky130_fd_sc_hd__and3_1
XFILLER_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08582_/C vssd1 vssd1 vccd1 vccd1 _08588_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _12418_/A vssd1 vssd1 vccd1 vccd1 _11560_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10511_ _10511_/A _10511_/B _10515_/B vssd1 vssd1 vccd1 vccd1 _15536_/D sky130_fd_sc_hd__nor3_1
XFILLER_128_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11491_ _11491_/A _11491_/B vssd1 vssd1 vccd1 vccd1 _11492_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13230_ _13281_/A _13230_/B _13230_/C vssd1 vssd1 vccd1 vccd1 _13231_/A sky130_fd_sc_hd__and3_1
X_10442_ _10439_/X _10440_/Y _10441_/Y _10437_/C vssd1 vssd1 vccd1 vccd1 _10444_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13161_ _15957_/Q _13193_/C _13041_/X vssd1 vssd1 vccd1 vccd1 _13163_/B sky130_fd_sc_hd__a21oi_1
X_10373_ _10663_/A vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12112_ _12112_/A _12112_/B _12112_/C vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__and3_1
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13092_ _13097_/C vssd1 vssd1 vccd1 vccd1 _13109_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12043_ _12039_/X _12040_/Y _12042_/Y _12037_/C vssd1 vssd1 vccd1 vccd1 _12045_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_123_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15802_ _07603_/A _15802_/D vssd1 vssd1 vccd1 vccd1 _15802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13994_ _14098_/A _13994_/B _13998_/B vssd1 vssd1 vccd1 vccd1 _16101_/D sky130_fd_sc_hd__nor3_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15733_ _15794_/CLK _15733_/D vssd1 vssd1 vccd1 vccd1 _15733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12945_ _12959_/A _12945_/B _12945_/C vssd1 vssd1 vccd1 vccd1 _12946_/A sky130_fd_sc_hd__and3_1
XFILLER_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15664_ _15763_/CLK _15664_/D vssd1 vssd1 vccd1 vccd1 _15664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12876_ _12896_/C vssd1 vssd1 vccd1 vccd1 _12908_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14615_ _13925_/X _14612_/B _14614_/X vssd1 vssd1 vccd1 vccd1 _14615_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _15744_/Q _11943_/B _11827_/C vssd1 vssd1 vccd1 vccd1 _11836_/A sky130_fd_sc_hd__and3_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _15194_/Q _15595_/D vssd1 vssd1 vccd1 vccd1 _15595_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11758_/A vssd1 vssd1 vccd1 vccd1 _15732_/D sky130_fd_sc_hd__clkbuf_1
X_14546_ _16219_/Q _14546_/B _14546_/C vssd1 vssd1 vccd1 vccd1 _14551_/A sky130_fd_sc_hd__and3_1
XFILLER_14_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10709_ _10710_/B _10710_/C _10710_/A vssd1 vssd1 vccd1 vccd1 _10711_/B sky130_fd_sc_hd__a21o_1
X_11689_ _15723_/Q _11863_/B _11689_/C vssd1 vssd1 vccd1 vccd1 _11689_/X sky130_fd_sc_hd__and3_1
X_14477_ _14471_/B _14472_/C _14481_/A _14475_/Y vssd1 vssd1 vccd1 vccd1 _14481_/B
+ sky130_fd_sc_hd__a211oi_1
X_16216_ _16240_/CLK _16216_/D vssd1 vssd1 vccd1 vccd1 _16216_/Q sky130_fd_sc_hd__dfxtp_2
X_13428_ _13481_/A _13428_/B _13428_/C vssd1 vssd1 vccd1 vccd1 _13429_/A sky130_fd_sc_hd__and3_1
X_16147_ _16148_/CLK _16147_/D vssd1 vssd1 vccd1 vccd1 _16147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13359_ _13358_/B _13358_/C _13305_/X vssd1 vssd1 vccd1 vccd1 _13360_/C sky130_fd_sc_hd__o21ai_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16078_ _16124_/CLK _16078_/D vssd1 vssd1 vccd1 vccd1 _16078_/Q sky130_fd_sc_hd__dfxtp_1
X_07920_ _07920_/A _07920_/B vssd1 vssd1 vccd1 vccd1 _07954_/B sky130_fd_sc_hd__xor2_4
X_15029_ _15029_/A vssd1 vssd1 vccd1 vccd1 _16325_/D sky130_fd_sc_hd__clkbuf_1
X_07851_ _15800_/Q vssd1 vssd1 vccd1 vccd1 _12193_/A sky130_fd_sc_hd__inv_2
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07782_ _15710_/Q _07783_/B vssd1 vssd1 vccd1 vccd1 _07784_/A sky130_fd_sc_hd__nand2_1
Xinput2 in1[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
X_09521_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09643_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09452_ _10896_/A vssd1 vssd1 vccd1 vccd1 _10610_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08403_ hold16/A _08403_/B vssd1 vssd1 vccd1 vccd1 _08415_/A sky130_fd_sc_hd__and2_1
X_09383_ _09377_/B _09378_/C _09380_/X _09381_/Y vssd1 vssd1 vccd1 vccd1 _09384_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08334_ _08722_/A vssd1 vssd1 vccd1 vccd1 _15086_/A sky130_fd_sc_hd__buf_4
XFILLER_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08265_ _08151_/A _08151_/B _08264_/Y vssd1 vssd1 vccd1 vccd1 _08266_/B sky130_fd_sc_hd__a21oi_2
X_08196_ _07979_/A _07979_/B _08195_/X vssd1 vssd1 vccd1 vccd1 _08287_/B sky130_fd_sc_hd__a21oi_2
XFILLER_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09719_ _15415_/Q _09950_/B _09727_/C vssd1 vssd1 vccd1 vccd1 _09724_/A sky130_fd_sc_hd__and3_1
XFILLER_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10991_ _11085_/A _10991_/B _10996_/A vssd1 vssd1 vccd1 vccd1 _15612_/D sky130_fd_sc_hd__nor3_1
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12727_/X _12728_/Y _12729_/Y _12724_/C vssd1 vssd1 vccd1 vccd1 _12732_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12661_/A vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__buf_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14400_ _14398_/A _14398_/B _14397_/Y _14399_/Y vssd1 vssd1 vccd1 vccd1 _16183_/D
+ sky130_fd_sc_hd__o31a_1
X_11612_ _11612_/A vssd1 vssd1 vccd1 vccd1 _11842_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _15484_/CLK _15380_/D vssd1 vssd1 vccd1 vccd1 _15380_/Q sky130_fd_sc_hd__dfxtp_1
X_12592_ _15865_/Q _12630_/C _12481_/X vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11543_ _15698_/Q _11601_/B _11547_/C vssd1 vssd1 vccd1 vccd1 _11543_/Y sky130_fd_sc_hd__nand3_1
X_14331_ _16187_/Q _16186_/Q _16185_/Q _14202_/X vssd1 vssd1 vccd1 vccd1 _16170_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14262_ _16159_/Q _14440_/B _14269_/C vssd1 vssd1 vccd1 vccd1 _14265_/A sky130_fd_sc_hd__and3_1
X_11474_ _15688_/Q _11650_/B _11479_/C vssd1 vssd1 vccd1 vccd1 _11474_/Y sky130_fd_sc_hd__nand3_1
XFILLER_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13213_ _13226_/C vssd1 vssd1 vccd1 vccd1 _13240_/C sky130_fd_sc_hd__clkbuf_1
X_16001_ _16011_/CLK _16001_/D vssd1 vssd1 vccd1 vccd1 _16001_/Q sky130_fd_sc_hd__dfxtp_2
X_10425_ _11634_/A vssd1 vssd1 vccd1 vccd1 _10654_/B sky130_fd_sc_hd__buf_2
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14193_ _14321_/A _14193_/B vssd1 vssd1 vccd1 vccd1 _14193_/Y sky130_fd_sc_hd__nor2_1
X_13144_ _13142_/A _13142_/B _13143_/X vssd1 vssd1 vccd1 vccd1 _15951_/D sky130_fd_sc_hd__a21oi_1
XFILLER_124_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10356_ _15515_/Q _10590_/B _10363_/C vssd1 vssd1 vccd1 vccd1 _10360_/B sky130_fd_sc_hd__nand3_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13075_ _13081_/A _13072_/Y _13074_/Y _13069_/C vssd1 vssd1 vccd1 vccd1 _13077_/B
+ sky130_fd_sc_hd__o211a_1
X_10287_ _10287_/A vssd1 vssd1 vccd1 vccd1 _15502_/D sky130_fd_sc_hd__clkbuf_1
X_12026_ _12084_/A _12026_/B _12030_/A vssd1 vssd1 vccd1 vccd1 _15774_/D sky130_fd_sc_hd__nor3_1
XFILLER_104_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13977_ _13990_/C vssd1 vssd1 vccd1 vccd1 _14003_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15716_ _15763_/CLK _15716_/D vssd1 vssd1 vccd1 vccd1 _15716_/Q sky130_fd_sc_hd__dfxtp_1
X_12928_ _15917_/Q vssd1 vssd1 vccd1 vccd1 _12941_/C sky130_fd_sc_hd__inv_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15647_ _15701_/CLK _15647_/D vssd1 vssd1 vccd1 vccd1 _15647_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12859_ _12857_/Y _12851_/C _12864_/A _12856_/Y vssd1 vssd1 vccd1 vccd1 _12864_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15578_ _15194_/Q _15578_/D vssd1 vssd1 vccd1 vccd1 _15578_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14529_ _14524_/Y _14527_/X _14528_/X vssd1 vssd1 vccd1 vccd1 _14529_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ _12249_/A _12361_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _08052_/C sky130_fd_sc_hd__o21a_1
XFILLER_128_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08952_ _15296_/Q _08951_/C _08888_/X vssd1 vssd1 vccd1 vccd1 _08953_/B sky130_fd_sc_hd__a21oi_1
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07903_ _13626_/C _07970_/B vssd1 vssd1 vccd1 vccd1 _07909_/A sky130_fd_sc_hd__xnor2_4
X_08883_ _08891_/A _08881_/Y _08882_/Y _08878_/C vssd1 vssd1 vccd1 vccd1 _08885_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07834_ _15836_/Q vssd1 vssd1 vccd1 vccd1 _12420_/A sky130_fd_sc_hd__clkinv_4
XFILLER_2_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07765_ _08099_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _07766_/B sky130_fd_sc_hd__xnor2_4
X_09504_ _15382_/Q _09733_/B _09508_/C vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__and3_1
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07696_ _13715_/A vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__buf_4
XFILLER_25_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09435_ _09435_/A _09435_/B _09435_/C vssd1 vssd1 vccd1 vccd1 _09436_/C sky130_fd_sc_hd__nand3_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09487_/A sky130_fd_sc_hd__buf_2
X_08317_ _08343_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _08359_/A sky130_fd_sc_hd__xnor2_2
X_09297_ _15350_/Q _09354_/B _09297_/C vssd1 vssd1 vccd1 vccd1 _09306_/B sky130_fd_sc_hd__and3_1
XANTENNA_40 _14892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _08249_/A _08249_/B _08249_/C vssd1 vssd1 vccd1 vccd1 _08250_/A sky130_fd_sc_hd__a21oi_1
XFILLER_138_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08179_ _08179_/A _08179_/B vssd1 vssd1 vccd1 vccd1 _08267_/A sky130_fd_sc_hd__nand2_2
X_10210_ _10210_/A _10210_/B _10210_/C vssd1 vssd1 vccd1 vccd1 _10211_/A sky130_fd_sc_hd__and3_1
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ _11190_/A vssd1 vssd1 vccd1 vccd1 _15643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10141_ _15481_/Q _10310_/B _10143_/C vssd1 vssd1 vccd1 vccd1 _10141_/X sky130_fd_sc_hd__and3_1
XFILLER_0_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10072_ _10097_/A _10072_/B _10072_/C vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__and3_1
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13900_ _13896_/A _13896_/B _13895_/Y _13899_/Y vssd1 vssd1 vccd1 vccd1 _16084_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14880_ _14880_/A _14880_/B vssd1 vssd1 vccd1 vccd1 _14881_/B sky130_fd_sc_hd__nor2_1
XFILLER_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13831_ _13831_/A vssd1 vssd1 vccd1 vccd1 _16073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10974_ _11551_/A vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__clkbuf_2
X_13762_ _14879_/A vssd1 vssd1 vccd1 vccd1 _14644_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15501_ _15224_/Q _15501_/D vssd1 vssd1 vccd1 vccd1 _15501_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12713_ _12713_/A vssd1 vssd1 vccd1 vccd1 _12935_/B sky130_fd_sc_hd__buf_2
X_13693_ _13693_/A vssd1 vssd1 vccd1 vccd1 _13693_/X sky130_fd_sc_hd__buf_2
X_15432_ _15483_/CLK _15432_/D vssd1 vssd1 vccd1 vccd1 _15432_/Q sky130_fd_sc_hd__dfxtp_2
X_12644_ _15880_/Q _15879_/Q _15878_/Q _12418_/X vssd1 vssd1 vccd1 vccd1 _15872_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15363_ _15377_/CLK _15363_/D vssd1 vssd1 vccd1 vccd1 _15363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12575_ _15862_/Q _12575_/B _12575_/C vssd1 vssd1 vccd1 vccd1 _12583_/B sky130_fd_sc_hd__and3_1
X_14314_ _16169_/Q _14313_/C _14270_/X vssd1 vssd1 vccd1 vccd1 _14315_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ _12100_/A vssd1 vssd1 vccd1 vccd1 _11526_/X sky130_fd_sc_hd__clkbuf_2
X_15294_ _15301_/CLK _15294_/D vssd1 vssd1 vccd1 vccd1 _15294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14245_ _14256_/C vssd1 vssd1 vccd1 vccd1 _14269_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11457_ _15687_/Q _11576_/B _11457_/C vssd1 vssd1 vccd1 vccd1 _11457_/X sky130_fd_sc_hd__and3_1
X_10408_ _10408_/A vssd1 vssd1 vccd1 vccd1 _15520_/D sky130_fd_sc_hd__clkbuf_1
X_14176_ _16141_/Q _14221_/B _14185_/C vssd1 vssd1 vccd1 vccd1 _14180_/A sky130_fd_sc_hd__and3_1
X_11388_ _11388_/A vssd1 vssd1 vccd1 vccd1 _11401_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10339_ _10337_/A _10337_/B _10338_/X vssd1 vssd1 vccd1 vccd1 _15510_/D sky130_fd_sc_hd__a21oi_1
X_13127_ _15952_/Q _14402_/A _13127_/C vssd1 vssd1 vccd1 vccd1 _13141_/A sky130_fd_sc_hd__and3_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _15941_/Q _13059_/C _13130_/A vssd1 vssd1 vccd1 vccd1 _13058_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12009_ _12015_/B _12009_/B vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__or2_1
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _13057_/B vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09151_ _09151_/A vssd1 vssd1 vccd1 vccd1 _15326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08102_ _08234_/A _08234_/B vssd1 vssd1 vccd1 vccd1 _08103_/B sky130_fd_sc_hd__xor2_4
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09202_/A sky130_fd_sc_hd__buf_2
X_08033_ _08033_/A _08033_/B _08033_/C vssd1 vssd1 vccd1 vccd1 _08034_/B sky130_fd_sc_hd__and3_1
XFILLER_128_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09984_ _09992_/A _09982_/Y _09983_/Y _09977_/C vssd1 vssd1 vccd1 vccd1 _09986_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08935_ _08935_/A vssd1 vssd1 vccd1 vccd1 _15292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08866_ _15284_/Q _08867_/C _08634_/X vssd1 vssd1 vccd1 vccd1 _08866_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07817_ _08052_/B _07817_/B vssd1 vssd1 vccd1 vccd1 _07818_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08797_ _15273_/Q _08802_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _08799_/C sky130_fd_sc_hd__a21o_1
XFILLER_84_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07748_ _15449_/Q _15431_/Q vssd1 vssd1 vccd1 vccd1 _07750_/A sky130_fd_sc_hd__or2_1
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ _07675_/X _07665_/A _07668_/B _07678_/Y vssd1 vssd1 vccd1 vccd1 _15202_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ _09536_/A vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__clkbuf_2
X_10690_ _10690_/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10694_/C sky130_fd_sc_hd__nor2_1
XFILLER_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09349_ _15358_/Q _09354_/C _09118_/X vssd1 vssd1 vccd1 vccd1 _09349_/Y sky130_fd_sc_hd__a21oi_1
X_12360_ _15835_/Q _15834_/Q _15833_/Q _12134_/X vssd1 vssd1 vccd1 vccd1 _15827_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ _15663_/Q _11367_/B _11311_/C vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__and3_1
XFILLER_148_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12291_ _15817_/Q _12291_/B _12291_/C vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__and3_1
XFILLER_4_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14030_ _14030_/A vssd1 vssd1 vccd1 vccd1 _16109_/D sky130_fd_sc_hd__clkbuf_1
X_11242_ _11249_/A _11242_/B _11242_/C vssd1 vssd1 vccd1 vccd1 _11243_/A sky130_fd_sc_hd__and3_1
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11173_ _11189_/A _11173_/B _11173_/C vssd1 vssd1 vccd1 vccd1 _11174_/A sky130_fd_sc_hd__and3_1
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10124_ _10155_/C vssd1 vssd1 vccd1 vccd1 _10162_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15981_ _15994_/CLK _15981_/D vssd1 vssd1 vccd1 vccd1 _15981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10055_ _10097_/A _10055_/B _10055_/C vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__and3_1
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14932_ _14932_/A _14932_/B vssd1 vssd1 vccd1 vccd1 _16303_/D sky130_fd_sc_hd__nor2_1
XFILLER_76_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14863_ _16293_/Q _14941_/B _14863_/C vssd1 vssd1 vccd1 vccd1 _14866_/B sky130_fd_sc_hd__nand3_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13814_ _13844_/A _13814_/B _13814_/C vssd1 vssd1 vccd1 vccd1 _13815_/A sky130_fd_sc_hd__and3_1
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14794_ _14993_/A vssd1 vssd1 vccd1 vccd1 _14953_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13745_ _16059_/Q _13752_/C _13693_/X vssd1 vssd1 vccd1 vccd1 _13745_/Y sky130_fd_sc_hd__a21oi_1
X_10957_ _15607_/Q _10963_/B _10957_/C vssd1 vssd1 vccd1 vccd1 _10957_/Y sky130_fd_sc_hd__nand3_1
XFILLER_73_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13676_ _13730_/A _13676_/B _13683_/A vssd1 vssd1 vccd1 vccd1 _16045_/D sky130_fd_sc_hd__nor3_1
X_10888_ _15598_/Q _10888_/B _10890_/C vssd1 vssd1 vccd1 vccd1 _10888_/X sky130_fd_sc_hd__and3_1
X_15415_ _15483_/CLK _15415_/D vssd1 vssd1 vccd1 vccd1 _15415_/Q sky130_fd_sc_hd__dfxtp_1
X_12627_ _12625_/Y _12621_/C _12634_/A _12624_/Y vssd1 vssd1 vccd1 vccd1 _12634_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_129_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15346_ _15348_/CLK _15346_/D vssd1 vssd1 vccd1 vccd1 _15346_/Q sky130_fd_sc_hd__dfxtp_1
X_12558_ _12558_/A vssd1 vssd1 vccd1 vccd1 _15858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ _11509_/A _11509_/B _11515_/A vssd1 vssd1 vccd1 vccd1 _15693_/D sky130_fd_sc_hd__nor3_1
X_15277_ _15286_/CLK _15277_/D vssd1 vssd1 vccd1 vccd1 _15277_/Q sky130_fd_sc_hd__dfxtp_1
X_12489_ _12510_/A _12489_/B _12489_/C vssd1 vssd1 vccd1 vccd1 _12490_/A sky130_fd_sc_hd__and3_1
X_14228_ _16151_/Q _14357_/B _14228_/C vssd1 vssd1 vccd1 vccd1 _14228_/X sky130_fd_sc_hd__and3_1
XFILLER_113_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _16138_/Q _14185_/C _14069_/X vssd1 vssd1 vccd1 vccd1 _14162_/B sky130_fd_sc_hd__a21oi_1
XFILLER_140_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08720_ _08893_/A _08724_/C vssd1 vssd1 vccd1 vccd1 _08720_/X sky130_fd_sc_hd__or2_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08651_ _15250_/Q _10963_/C _08651_/C vssd1 vssd1 vccd1 vccd1 _08660_/A sky130_fd_sc_hd__and3_1
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07602_ _15195_/Q _08471_/B vssd1 vssd1 vccd1 vccd1 _15195_/D sky130_fd_sc_hd__nor2_1
XFILLER_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08582_ _15241_/Q _10963_/C _08582_/C vssd1 vssd1 vccd1 vccd1 _08593_/A sky130_fd_sc_hd__and3_1
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ _10065_/A vssd1 vssd1 vccd1 vccd1 _09432_/B sky130_fd_sc_hd__buf_2
XFILLER_148_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09134_ _09133_/B _09133_/C _09019_/X vssd1 vssd1 vccd1 vccd1 _09135_/C sky130_fd_sc_hd__o21ai_1
XFILLER_148_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09065_ _09063_/Y _09058_/C _09070_/A _09062_/Y vssd1 vssd1 vccd1 vccd1 _09070_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_147_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08016_ _08016_/A _07883_/B vssd1 vssd1 vccd1 vccd1 _08016_/X sky130_fd_sc_hd__or2b_1
XFILLER_118_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09967_ _15453_/Q _10199_/B _09967_/C vssd1 vssd1 vccd1 vccd1 _09967_/Y sky130_fd_sc_hd__nand3_1
XFILLER_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08918_ _08918_/A vssd1 vssd1 vccd1 vccd1 _15290_/D sky130_fd_sc_hd__clkbuf_1
X_09898_ _15443_/Q _09903_/C _09778_/X vssd1 vssd1 vccd1 vccd1 _09900_/C sky130_fd_sc_hd__a21o_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ input1/X vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__buf_6
XFILLER_85_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11860_ _11860_/A _11860_/B _11860_/C vssd1 vssd1 vccd1 vccd1 _11861_/C sky130_fd_sc_hd__nand3_1
XFILLER_73_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ _11099_/A vssd1 vssd1 vccd1 vccd1 _10931_/A sky130_fd_sc_hd__buf_2
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11791_ _11814_/C vssd1 vssd1 vccd1 vccd1 _11827_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_41_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ _13538_/A _13530_/B _13530_/C vssd1 vssd1 vccd1 vccd1 _13531_/A sky130_fd_sc_hd__and3_1
X_10742_ _15574_/Q _10741_/C _10624_/X vssd1 vssd1 vccd1 vccd1 _10743_/B sky130_fd_sc_hd__a21oi_1
XFILLER_25_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10673_ _15562_/Q _10729_/B _10679_/C vssd1 vssd1 vccd1 vccd1 _10673_/Y sky130_fd_sc_hd__nand3_1
XFILLER_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13461_ _13460_/B _13460_/C _13305_/X vssd1 vssd1 vccd1 vccd1 _13462_/C sky130_fd_sc_hd__o21ai_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15200_ _16359_/CLK _15200_/D vssd1 vssd1 vccd1 vccd1 _15200_/Q sky130_fd_sc_hd__dfxtp_2
X_12412_ _12410_/A _12410_/B _12411_/X vssd1 vssd1 vccd1 vccd1 _15834_/D sky130_fd_sc_hd__a21oi_1
X_16180_ _16189_/CLK _16180_/D vssd1 vssd1 vccd1 vccd1 _16180_/Q sky130_fd_sc_hd__dfxtp_2
X_13392_ _13410_/A _13392_/B _13392_/C vssd1 vssd1 vccd1 vccd1 _13393_/A sky130_fd_sc_hd__and3_1
X_15131_ _16356_/Q _15131_/B _15131_/C vssd1 vssd1 vccd1 vccd1 _15134_/B sky130_fd_sc_hd__nand3_1
X_12343_ _12341_/Y _12337_/C _12350_/A _12340_/Y vssd1 vssd1 vccd1 vccd1 _12350_/B
+ sky130_fd_sc_hd__a211oi_1
X_15062_ hold21/A _15061_/C _14942_/X vssd1 vssd1 vccd1 vccd1 _15064_/C sky130_fd_sc_hd__a21o_1
X_12274_ _12274_/A vssd1 vssd1 vccd1 vccd1 _15813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11225_ _11225_/A _11225_/B _11225_/C vssd1 vssd1 vccd1 vccd1 _11226_/C sky130_fd_sc_hd__nand3_1
X_14013_ _13921_/X _14011_/B _13922_/X vssd1 vssd1 vccd1 vccd1 _14013_/Y sky130_fd_sc_hd__a21oi_1
X_11156_ _11156_/A vssd1 vssd1 vccd1 vccd1 _11169_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10107_ _15475_/Q _10106_/C _10044_/X vssd1 vssd1 vccd1 vccd1 _10108_/B sky130_fd_sc_hd__a21oi_1
X_11087_ _15628_/Q _11086_/C _10911_/X vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__a21oi_1
X_15964_ _15970_/CLK _15964_/D vssd1 vssd1 vccd1 vccd1 _15964_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10038_ _15465_/Q _10043_/C _09981_/X vssd1 vssd1 vccd1 vccd1 _10038_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14915_ _14915_/A _14915_/B _14920_/B vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__nor3_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15895_ _07603_/A _15895_/D vssd1 vssd1 vccd1 vccd1 _15895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14846_ _14840_/A _14843_/B _14845_/X vssd1 vssd1 vccd1 vccd1 _14853_/C sky130_fd_sc_hd__o21a_1
XFILLER_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14777_ _16274_/Q _14795_/C _14702_/X vssd1 vssd1 vccd1 vccd1 _14779_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11989_ _11997_/A _11989_/B _11989_/C vssd1 vssd1 vccd1 vccd1 _11990_/A sky130_fd_sc_hd__and3_1
X_13728_ _16056_/Q _13758_/C _13573_/X vssd1 vssd1 vccd1 vccd1 _13730_/B sky130_fd_sc_hd__a21oi_1
X_13659_ _13659_/A _13659_/B vssd1 vssd1 vccd1 vccd1 _13662_/C sky130_fd_sc_hd__nor2_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15329_ _15337_/CLK _15329_/D vssd1 vssd1 vccd1 vccd1 _15329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09821_ _10110_/A vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09752_ _09750_/Y _09746_/C _09758_/A _09749_/Y vssd1 vssd1 vccd1 vccd1 _09758_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08703_ _08701_/Y _08697_/C _08699_/X _08700_/Y vssd1 vssd1 vccd1 vccd1 _08704_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09683_ _09690_/A _09683_/B _09683_/C vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__and3_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _13057_/B vssd1 vssd1 vccd1 vccd1 _08634_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08565_/A vssd1 vssd1 vccd1 vccd1 _15237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08496_ _08488_/B _08489_/C _08493_/X _08494_/Y vssd1 vssd1 vccd1 vccd1 _08497_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09117_ _15322_/Q _09290_/B _09117_/C vssd1 vssd1 vccd1 vccd1 _09128_/A sky130_fd_sc_hd__and3_1
XFILLER_148_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09048_ _09045_/X _09046_/Y _09047_/Y _09043_/C vssd1 vssd1 vccd1 vccd1 _09050_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_124_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _11008_/Y _11003_/C _11006_/X _11007_/Y vssd1 vssd1 vccd1 vccd1 _11011_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12961_ _13239_/A vssd1 vssd1 vccd1 vccd1 _13077_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14700_ _16268_/Q _16267_/Q _16266_/Q _14620_/X vssd1 vssd1 vccd1 vccd1 _16251_/D
+ sky130_fd_sc_hd__o31a_1
X_11912_ _13041_/A vssd1 vssd1 vccd1 vccd1 _11912_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _15763_/CLK _15680_/D vssd1 vssd1 vccd1 vccd1 _15680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _12892_/A vssd1 vssd1 vccd1 vccd1 _15911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14748_/A _14631_/B _14631_/C vssd1 vssd1 vccd1 vccd1 _14632_/A sky130_fd_sc_hd__and3_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11843_ _12015_/A _11843_/B _11843_/C vssd1 vssd1 vccd1 vccd1 _11845_/B sky130_fd_sc_hd__or3_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _14562_/A _14562_/B vssd1 vssd1 vccd1 vccd1 _14562_/X sky130_fd_sc_hd__or2_1
X_11774_ _15736_/Q _12007_/B _11774_/C vssd1 vssd1 vccd1 vccd1 _11784_/B sky130_fd_sc_hd__and3_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16312_/CLK _16301_/D vssd1 vssd1 vccd1 vccd1 _16301_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13512_/B _13512_/C _13305_/X vssd1 vssd1 vccd1 vccd1 _13514_/C sky130_fd_sc_hd__o21ai_1
X_10725_ _10732_/A _10725_/B _10725_/C vssd1 vssd1 vccd1 vccd1 _10726_/A sky130_fd_sc_hd__and3_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _14533_/A _14493_/B vssd1 vssd1 vccd1 vccd1 _14493_/Y sky130_fd_sc_hd__nor2_1
X_16232_ _16367_/CLK _16232_/D vssd1 vssd1 vccd1 vccd1 _16232_/Q sky130_fd_sc_hd__dfxtp_1
X_13444_ _13700_/A vssd1 vssd1 vccd1 vccd1 _13648_/B sky130_fd_sc_hd__clkbuf_4
X_10656_ _15561_/Q _10665_/C _10655_/X vssd1 vssd1 vccd1 vccd1 _10656_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16163_ _16187_/CLK _16163_/D vssd1 vssd1 vccd1 vccd1 _16163_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10587_ _11507_/A vssd1 vssd1 vccd1 vccd1 _10817_/B sky130_fd_sc_hd__clkbuf_4
X_13375_ _15994_/Q _13380_/C _13269_/X vssd1 vssd1 vccd1 vccd1 _13377_/C sky130_fd_sc_hd__a21o_1
X_15114_ _15109_/A _15112_/B _15043_/X vssd1 vssd1 vccd1 vccd1 _15120_/C sky130_fd_sc_hd__o21a_1
X_12326_ _15822_/Q _12554_/B _12326_/C vssd1 vssd1 vccd1 vccd1 _12326_/Y sky130_fd_sc_hd__nand3_1
XFILLER_126_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16094_ _16224_/CLK _16094_/D vssd1 vssd1 vccd1 vccd1 _16094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15045_ _15045_/A _15051_/C vssd1 vssd1 vccd1 vccd1 _15045_/Y sky130_fd_sc_hd__nor2_1
X_12257_ _15812_/Q _12262_/C _12086_/X vssd1 vssd1 vccd1 vccd1 _12259_/C sky130_fd_sc_hd__a21o_1
XFILLER_141_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11208_ _11439_/A _11208_/B _11208_/C vssd1 vssd1 vccd1 vccd1 _11210_/B sky130_fd_sc_hd__or3_1
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12188_ _12188_/A vssd1 vssd1 vccd1 vccd1 _12188_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _15635_/Q _11313_/B _11143_/C vssd1 vssd1 vccd1 vccd1 _11139_/Y sky130_fd_sc_hd__nand3_1
X_15947_ _16100_/CLK _15947_/D vssd1 vssd1 vccd1 vccd1 _15947_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15878_ _15907_/CLK _15878_/D vssd1 vssd1 vccd1 vccd1 _15878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14829_ _14829_/A _14829_/B _14829_/C vssd1 vssd1 vccd1 vccd1 _14830_/C sky130_fd_sc_hd__nand3_1
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08350_ _08386_/B _08350_/B vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__and2_1
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08281_ _08272_/A _08272_/B _08271_/A vssd1 vssd1 vccd1 vccd1 _08330_/A sky130_fd_sc_hd__a21oi_2
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09804_ _15427_/Q _09862_/B _09811_/C vssd1 vssd1 vccd1 vccd1 _09804_/Y sky130_fd_sc_hd__nand3_1
XFILLER_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07996_ _16161_/Q _07996_/B vssd1 vssd1 vccd1 vccd1 _07996_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09735_ _15417_/Q _09911_/B _09735_/C vssd1 vssd1 vccd1 vccd1 _09735_/Y sky130_fd_sc_hd__nand3_1
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09666_ _15407_/Q _09671_/C _09490_/X vssd1 vssd1 vccd1 vccd1 _09668_/C sky130_fd_sc_hd__a21o_1
XFILLER_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _15246_/Q _08622_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _08619_/C sky130_fd_sc_hd__a21o_1
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09594_/B _09594_/C _09596_/X vssd1 vssd1 vccd1 vccd1 _09598_/C sky130_fd_sc_hd__o21ai_1
XFILLER_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08568_/C vssd1 vssd1 vccd1 vccd1 _08582_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08479_ input1/X vssd1 vssd1 vccd1 vccd1 _12650_/A sky130_fd_sc_hd__buf_4
X_10510_ _10508_/Y _10503_/C _10515_/A _10507_/Y vssd1 vssd1 vccd1 vccd1 _10515_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11490_ _11497_/B _11490_/B vssd1 vssd1 vccd1 vccd1 _11492_/A sky130_fd_sc_hd__or2_1
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ _15526_/Q _10441_/B _10446_/C vssd1 vssd1 vccd1 vccd1 _10441_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10372_ _15517_/Q _10602_/B _10375_/C vssd1 vssd1 vccd1 vccd1 _10372_/X sky130_fd_sc_hd__and3_1
X_13160_ _13187_/C vssd1 vssd1 vccd1 vccd1 _13193_/C sky130_fd_sc_hd__clkbuf_2
X_12111_ _12109_/Y _12105_/C _12107_/X _12108_/Y vssd1 vssd1 vccd1 vccd1 _12112_/C
+ sky130_fd_sc_hd__a211o_1
X_13091_ _13239_/A vssd1 vssd1 vccd1 vccd1 _13218_/A sky130_fd_sc_hd__buf_2
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12042_ _15777_/Q _12270_/B _12042_/C vssd1 vssd1 vccd1 vccd1 _12042_/Y sky130_fd_sc_hd__nand3_1
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15801_ _07603_/A _15801_/D vssd1 vssd1 vccd1 vccd1 _15801_/Q sky130_fd_sc_hd__dfxtp_2
X_13993_ _13985_/B _13986_/C _13998_/A _13991_/Y vssd1 vssd1 vccd1 vccd1 _13998_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15732_ _15794_/CLK _15732_/D vssd1 vssd1 vccd1 vccd1 _15732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _12938_/B _12939_/C _12941_/X _12942_/Y vssd1 vssd1 vccd1 vccd1 _12945_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_73_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15663_ _15763_/CLK _15663_/D vssd1 vssd1 vccd1 vccd1 _15663_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12875_ _12887_/C vssd1 vssd1 vccd1 vccd1 _12896_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _15014_/A vssd1 vssd1 vccd1 vccd1 _14614_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _11826_/A vssd1 vssd1 vccd1 vccd1 _11949_/A sky130_fd_sc_hd__buf_2
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15194_/Q _15594_/D vssd1 vssd1 vccd1 vccd1 _15594_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _16219_/Q _14566_/C _14503_/X vssd1 vssd1 vccd1 vccd1 _14547_/B sky130_fd_sc_hd__a21oi_1
X_11757_ _11765_/A _11757_/B _11757_/C vssd1 vssd1 vccd1 vccd1 _11758_/A sky130_fd_sc_hd__and3_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ _15569_/Q _10714_/C _10648_/X vssd1 vssd1 vccd1 vccd1 _10710_/C sky130_fd_sc_hd__a21o_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14476_ _14481_/A _14475_/Y _14471_/B _14472_/C vssd1 vssd1 vccd1 vccd1 _14478_/B
+ sky130_fd_sc_hd__o211a_1
X_11688_ _11688_/A vssd1 vssd1 vccd1 vccd1 _15721_/D sky130_fd_sc_hd__clkbuf_1
X_16215_ _16367_/CLK _16215_/D vssd1 vssd1 vccd1 vccd1 _16215_/Q sky130_fd_sc_hd__dfxtp_2
X_13427_ _13427_/A _13427_/B _13427_/C vssd1 vssd1 vccd1 vccd1 _13428_/C sky130_fd_sc_hd__nand3_1
X_10639_ _10639_/A vssd1 vssd1 vccd1 vccd1 _10654_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16146_ _16166_/CLK _16146_/D vssd1 vssd1 vccd1 vccd1 _16146_/Q sky130_fd_sc_hd__dfxtp_2
X_13358_ _13408_/A _13358_/B _13358_/C vssd1 vssd1 vccd1 vccd1 _13360_/B sky130_fd_sc_hd__or3_1
X_12309_ _15820_/Q _12309_/B _12317_/C vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__and3_1
X_16077_ _16124_/CLK _16077_/D vssd1 vssd1 vccd1 vccd1 _16077_/Q sky130_fd_sc_hd__dfxtp_1
X_13289_ _13339_/A _13289_/B _13289_/C vssd1 vssd1 vccd1 vccd1 _13290_/A sky130_fd_sc_hd__and3_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15028_ _15135_/A _15028_/B _15028_/C vssd1 vssd1 vccd1 vccd1 _15029_/A sky130_fd_sc_hd__and3_1
XFILLER_114_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07850_ _15782_/Q vssd1 vssd1 vccd1 vccd1 _12077_/A sky130_fd_sc_hd__clkinv_4
XFILLER_110_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07781_ _08083_/A _07781_/B vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__xnor2_1
Xinput3 in1[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
X_09520_ _09520_/A vssd1 vssd1 vccd1 vccd1 _15382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09451_ _15374_/Q _09451_/B _09460_/C vssd1 vssd1 vccd1 vccd1 _09451_/X sky130_fd_sc_hd__and3_1
X_08402_ _08375_/A _08375_/B _08397_/B _08397_/A _08372_/A vssd1 vssd1 vccd1 vccd1
+ _08411_/C sky130_fd_sc_hd__o221a_1
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09382_ _09380_/X _09381_/Y _09377_/B _09378_/C vssd1 vssd1 vccd1 vccd1 _09384_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_52_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ _08274_/Y _08276_/Y _08332_/Y vssd1 vssd1 vccd1 vccd1 _08333_/X sky130_fd_sc_hd__o21a_1
X_08264_ _08264_/A _08264_/B vssd1 vssd1 vccd1 vccd1 _08264_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08195_ _07978_/B _08195_/B vssd1 vssd1 vccd1 vccd1 _08195_/X sky130_fd_sc_hd__and2b_1
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07979_ _07979_/A _07979_/B vssd1 vssd1 vccd1 vccd1 _08180_/A sky130_fd_sc_hd__xnor2_2
X_09718_ _10007_/A vssd1 vssd1 vccd1 vccd1 _09950_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10990_ _15613_/Q _11161_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _10996_/A sky130_fd_sc_hd__and3_1
XFILLER_16_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09649_ _09760_/A _09652_/C vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__or2_1
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _15876_/Q _12720_/B _12660_/C vssd1 vssd1 vccd1 vccd1 _12660_/X sky130_fd_sc_hd__and3_1
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11609_/A _11609_/B _11610_/X vssd1 vssd1 vccd1 vccd1 _15708_/D sky130_fd_sc_hd__a21oi_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12591_ _12623_/C vssd1 vssd1 vccd1 vccd1 _12630_/C sky130_fd_sc_hd__clkbuf_2
X_14330_ _14330_/A _14330_/B vssd1 vssd1 vccd1 vccd1 _16169_/D sky130_fd_sc_hd__nor2_1
X_11542_ _15699_/Q _11547_/C _11425_/X vssd1 vssd1 vccd1 vccd1 _11542_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14261_ _14261_/A vssd1 vssd1 vccd1 vccd1 _14440_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11473_ _15689_/Q _11479_/C _11472_/X vssd1 vssd1 vccd1 vccd1 _11473_/Y sky130_fd_sc_hd__a21oi_1
X_16000_ _16007_/CLK _16000_/D vssd1 vssd1 vccd1 vccd1 _16000_/Q sky130_fd_sc_hd__dfxtp_2
X_13212_ _13217_/C vssd1 vssd1 vccd1 vccd1 _13226_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10424_ input3/X vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__buf_2
X_14192_ _14320_/A _14192_/B vssd1 vssd1 vccd1 vccd1 _14193_/B sky130_fd_sc_hd__and2_1
XFILLER_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13143_ _13199_/A _13146_/C vssd1 vssd1 vccd1 vccd1 _13143_/X sky130_fd_sc_hd__or2_1
X_10355_ _11569_/A vssd1 vssd1 vccd1 vccd1 _10590_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10323_/A _10286_/B _10286_/C vssd1 vssd1 vccd1 vccd1 _10287_/A sky130_fd_sc_hd__and3_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _15942_/Q _14402_/A _13078_/C vssd1 vssd1 vccd1 vccd1 _13074_/Y sky130_fd_sc_hd__nand3_1
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12025_ _15775_/Q _12025_/B _12033_/C vssd1 vssd1 vccd1 vccd1 _12030_/A sky130_fd_sc_hd__and3_1
XFILLER_116_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13976_ _13979_/C vssd1 vssd1 vccd1 vccd1 _13990_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15715_ _15794_/CLK _15715_/D vssd1 vssd1 vccd1 vccd1 _15715_/Q sky130_fd_sc_hd__dfxtp_1
X_12927_ _15923_/Q _15925_/Q _15924_/Q _12704_/X vssd1 vssd1 vccd1 vccd1 _15917_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15646_ _15655_/CLK _15646_/D vssd1 vssd1 vccd1 vccd1 _15646_/Q sky130_fd_sc_hd__dfxtp_1
X_12858_ _12864_/A _12856_/Y _12857_/Y _12851_/C vssd1 vssd1 vccd1 vccd1 _12860_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ _11824_/A _11809_/B _11809_/C vssd1 vssd1 vccd1 vccd1 _11810_/A sky130_fd_sc_hd__and3_1
XFILLER_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15577_ _15194_/Q _15577_/D vssd1 vssd1 vccd1 vccd1 _15577_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12796_/A _12789_/B _12789_/C vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__and3_1
XFILLER_42_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14528_ _15014_/A vssd1 vssd1 vccd1 vccd1 _14528_/X sky130_fd_sc_hd__clkbuf_2
X_14459_ _14459_/A vssd1 vssd1 vccd1 vccd1 _14459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16129_ _16129_/CLK _16129_/D vssd1 vssd1 vccd1 vccd1 _16129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08951_ _15296_/Q _09067_/B _08951_/C vssd1 vssd1 vccd1 vccd1 _08961_/B sky130_fd_sc_hd__and3_1
XFILLER_142_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07902_ _16215_/Q _07967_/B vssd1 vssd1 vccd1 vccd1 _07970_/B sky130_fd_sc_hd__xnor2_4
X_08882_ _15285_/Q _08947_/B _08886_/C vssd1 vssd1 vccd1 vccd1 _08882_/Y sky130_fd_sc_hd__nand3_1
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07833_ _15656_/Q vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__clkinv_2
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07764_ _15521_/Q _08093_/B vssd1 vssd1 vccd1 vccd1 _08100_/B sky130_fd_sc_hd__xnor2_4
XFILLER_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09503_ _10081_/A vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__buf_2
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07695_ _12631_/A vssd1 vssd1 vccd1 vccd1 _13715_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09434_ _09435_/B _09435_/C _09435_/A vssd1 vssd1 vccd1 vccd1 _09436_/B sky130_fd_sc_hd__a21o_1
XFILLER_25_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _09365_/A vssd1 vssd1 vccd1 vccd1 _15359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08316_ _08349_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__and2_1
X_09296_ _09353_/A _09296_/B _09300_/B vssd1 vssd1 vccd1 vccd1 _15348_/D sky130_fd_sc_hd__nor3_1
XANTENNA_30 _14892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08247_ _08131_/A _08131_/B _08384_/A _08246_/X vssd1 vssd1 vccd1 vccd1 _08249_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08178_ _08178_/A _07985_/B vssd1 vssd1 vccd1 vccd1 _08179_/B sky130_fd_sc_hd__or2b_1
XFILLER_134_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10140_ _10140_/A vssd1 vssd1 vccd1 vccd1 _15479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10071_ _10071_/A _10071_/B _10071_/C vssd1 vssd1 vccd1 vccd1 _10072_/C sky130_fd_sc_hd__nand3_1
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13830_ _13844_/A _13830_/B _13830_/C vssd1 vssd1 vccd1 vccd1 _13831_/A sky130_fd_sc_hd__and3_1
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ _13761_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13763_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10973_ _10973_/A _10973_/B vssd1 vssd1 vccd1 vccd1 _10975_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15500_ _15224_/Q _15500_/D vssd1 vssd1 vccd1 vccd1 _15500_/Q sky130_fd_sc_hd__dfxtp_1
X_12712_ _12804_/A _12712_/B _12717_/A vssd1 vssd1 vccd1 vccd1 _15882_/D sky130_fd_sc_hd__nor3_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _16050_/Q _13838_/B _13701_/C vssd1 vssd1 vccd1 vccd1 _13692_/X sky130_fd_sc_hd__and3_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15431_ _15440_/CLK _15431_/D vssd1 vssd1 vccd1 vccd1 _15431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12643_ _12643_/A vssd1 vssd1 vccd1 vccd1 _15871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ _15377_/CLK _15362_/D vssd1 vssd1 vccd1 vccd1 _15362_/Q sky130_fd_sc_hd__dfxtp_1
X_12574_ _12652_/A _12574_/B _12578_/B vssd1 vssd1 vccd1 vccd1 _15860_/D sky130_fd_sc_hd__nor3_1
XFILLER_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14313_ _16169_/Q _14357_/B _14313_/C vssd1 vssd1 vccd1 vccd1 _14313_/X sky130_fd_sc_hd__and3_1
X_11525_ _15697_/Q _11525_/B _11528_/C vssd1 vssd1 vccd1 vccd1 _11525_/X sky130_fd_sc_hd__and3_1
X_15293_ _15301_/CLK _15293_/D vssd1 vssd1 vccd1 vccd1 _15293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14244_ _14247_/C vssd1 vssd1 vccd1 vccd1 _14256_/C sky130_fd_sc_hd__clkbuf_1
X_11456_ _11456_/A vssd1 vssd1 vccd1 vccd1 _15685_/D sky130_fd_sc_hd__clkbuf_1
X_10407_ _10444_/A _10407_/B _10407_/C vssd1 vssd1 vccd1 vccd1 _10408_/A sky130_fd_sc_hd__and3_1
XFILLER_109_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14175_ _14208_/A _14175_/B _14179_/B vssd1 vssd1 vccd1 vccd1 _16137_/D sky130_fd_sc_hd__nor3_1
X_11387_ _11826_/A vssd1 vssd1 vccd1 vccd1 _11509_/A sky130_fd_sc_hd__buf_2
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13126_ _13126_/A vssd1 vssd1 vccd1 vccd1 _15949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10338_ _10338_/A _10342_/C vssd1 vssd1 vccd1 vccd1 _10338_/X sky130_fd_sc_hd__or2_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _15941_/Q _13057_/B _13059_/C vssd1 vssd1 vccd1 vccd1 _13057_/X sky130_fd_sc_hd__and3_1
X_10269_ _11137_/A vssd1 vssd1 vccd1 vccd1 _10269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12008_ _15772_/Q _12007_/C _11775_/X vssd1 vssd1 vccd1 vccd1 _12009_/B sky130_fd_sc_hd__a21oi_1
XFILLER_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13959_ _13957_/X _13959_/B vssd1 vssd1 vccd1 vccd1 _13959_/X sky130_fd_sc_hd__and2b_1
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15629_ _15665_/CLK _15629_/D vssd1 vssd1 vccd1 vccd1 _15629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09150_ _09171_/A _09150_/B _09150_/C vssd1 vssd1 vccd1 vccd1 _09151_/A sky130_fd_sc_hd__and3_1
XFILLER_147_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08101_ _14782_/C _07766_/B _08100_/X vssd1 vssd1 vccd1 vccd1 _08234_/B sky130_fd_sc_hd__o21a_4
X_09081_ _11963_/A vssd1 vssd1 vccd1 vccd1 _09657_/A sky130_fd_sc_hd__clkbuf_4
X_08032_ _08033_/A _08033_/B _08033_/C vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__a21oi_2
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ _15455_/Q _10102_/B _09989_/C vssd1 vssd1 vccd1 vccd1 _09983_/Y sky130_fd_sc_hd__nand3_1
XFILLER_115_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08934_ _08942_/A _08934_/B _08934_/C vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__and3_1
XFILLER_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08865_ _15284_/Q _08865_/B _08867_/C vssd1 vssd1 vccd1 vccd1 _08865_/X sky130_fd_sc_hd__and3_1
XFILLER_84_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07816_ _08052_/A _07815_/C _15791_/Q vssd1 vssd1 vccd1 vccd1 _07817_/B sky130_fd_sc_hd__a21o_1
X_08796_ _15273_/Q _08853_/B _08802_/C vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__nand3_1
XFILLER_38_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07747_ _15467_/Q vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__inv_2
XFILLER_38_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07678_ _14648_/A _07698_/C vssd1 vssd1 vccd1 vccd1 _07678_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09417_ _09415_/A _09415_/B _09416_/X vssd1 vssd1 vccd1 vccd1 _15366_/D sky130_fd_sc_hd__a21oi_1
XFILLER_13_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09348_ _15358_/Q _09577_/B _09348_/C vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__and3_1
XFILLER_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _09276_/X _09277_/Y _09278_/Y _09274_/C vssd1 vssd1 vccd1 vccd1 _09281_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _11310_/A vssd1 vssd1 vccd1 vccd1 _15661_/D sky130_fd_sc_hd__clkbuf_1
X_12290_ _12368_/A _12290_/B _12294_/B vssd1 vssd1 vccd1 vccd1 _15815_/D sky130_fd_sc_hd__nor3_1
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ _11239_/Y _11234_/C _11236_/X _11238_/Y vssd1 vssd1 vccd1 vccd1 _11242_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11172_ _11166_/B _11167_/C _11169_/X _11170_/Y vssd1 vssd1 vccd1 vccd1 _11173_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10123_ _10143_/C vssd1 vssd1 vccd1 vccd1 _10155_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15980_ _15984_/CLK _15980_/D vssd1 vssd1 vccd1 vccd1 _15980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ _10053_/B _10053_/C _09884_/X vssd1 vssd1 vccd1 vccd1 _10055_/C sky130_fd_sc_hd__o21ai_1
X_14931_ _14892_/X _14929_/A _14893_/X vssd1 vssd1 vccd1 vccd1 _14932_/B sky130_fd_sc_hd__o21ai_1
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14862_ _14915_/A _14862_/B _14866_/A vssd1 vssd1 vccd1 vccd1 _16288_/D sky130_fd_sc_hd__nor3_1
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13813_ _13812_/B _13812_/C _13919_/A vssd1 vssd1 vccd1 vccd1 _13814_/C sky130_fd_sc_hd__o21ai_1
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14793_ _14825_/A _14793_/B _14798_/B vssd1 vssd1 vccd1 vccd1 _16272_/D sky130_fd_sc_hd__nor3_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13744_ _16059_/Q _13838_/B _13752_/C vssd1 vssd1 vccd1 vccd1 _13744_/X sky130_fd_sc_hd__and3_1
X_10956_ _15608_/Q _10963_/B _10897_/X vssd1 vssd1 vccd1 vccd1 _10956_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13675_ _16047_/Q _13675_/B _13675_/C vssd1 vssd1 vccd1 vccd1 _13683_/A sky130_fd_sc_hd__and3_1
XFILLER_71_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10887_ _10887_/A vssd1 vssd1 vccd1 vccd1 _15596_/D sky130_fd_sc_hd__clkbuf_1
X_15414_ _15483_/CLK _15414_/D vssd1 vssd1 vccd1 vccd1 _15414_/Q sky130_fd_sc_hd__dfxtp_2
X_12626_ _12634_/A _12624_/Y _12625_/Y _12621_/C vssd1 vssd1 vccd1 vccd1 _12628_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15345_ _15348_/CLK _15345_/D vssd1 vssd1 vccd1 vccd1 _15345_/Q sky130_fd_sc_hd__dfxtp_1
X_12557_ _12565_/A _12557_/B _12557_/C vssd1 vssd1 vccd1 vccd1 _12558_/A sky130_fd_sc_hd__and3_1
XFILLER_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11508_ _15694_/Q _11737_/B _11518_/C vssd1 vssd1 vccd1 vccd1 _11515_/A sky130_fd_sc_hd__and3_1
X_15276_ _15286_/CLK _15276_/D vssd1 vssd1 vccd1 vccd1 _15276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12488_ _12488_/A _12488_/B _12488_/C vssd1 vssd1 vccd1 vccd1 _12489_/C sky130_fd_sc_hd__nand3_1
X_14227_ _14224_/B _14223_/Y _14224_/A vssd1 vssd1 vccd1 vccd1 _14227_/Y sky130_fd_sc_hd__o21bai_1
X_11439_ _11439_/A _11439_/B _11439_/C vssd1 vssd1 vccd1 vccd1 _11441_/B sky130_fd_sc_hd__or3_1
XFILLER_98_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14158_ _14171_/C vssd1 vssd1 vccd1 vccd1 _14185_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _15950_/Q _14298_/A _13109_/C vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__and3_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14089_ _14086_/X _14087_/Y _14088_/Y _14084_/C vssd1 vssd1 vccd1 vccd1 _14091_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08650_ _08944_/A vssd1 vssd1 vccd1 vccd1 _08774_/A sky130_fd_sc_hd__buf_2
XFILLER_94_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07601_ _15194_/Q _08471_/B vssd1 vssd1 vccd1 vccd1 _15194_/D sky130_fd_sc_hd__nor2_1
XFILLER_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08581_ _08581_/A vssd1 vssd1 vccd1 vccd1 _15239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09202_ _09202_/A _09202_/B _09208_/A vssd1 vssd1 vccd1 vccd1 _15334_/D sky130_fd_sc_hd__nor3_1
XFILLER_50_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09133_ _09133_/A _09133_/B _09133_/C vssd1 vssd1 vccd1 vccd1 _09135_/B sky130_fd_sc_hd__or3_1
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09064_ _09070_/A _09062_/Y _09063_/Y _09058_/C vssd1 vssd1 vccd1 vccd1 _09066_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08015_ _08205_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08019_/A sky130_fd_sc_hd__xnor2_1
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09966_ _10548_/A vssd1 vssd1 vccd1 vccd1 _10199_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_58_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08917_ _08942_/A _08917_/B _08917_/C vssd1 vssd1 vccd1 vccd1 _08918_/A sky130_fd_sc_hd__and3_1
XFILLER_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09897_ _15443_/Q _10010_/B _09903_/C vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__nand3_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08848_ _15281_/Q _08886_/C _08735_/X vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__a21oi_1
XFILLER_18_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08779_ _08779_/A _08779_/B vssd1 vssd1 vccd1 vccd1 _08783_/C sky130_fd_sc_hd__nor2_1
XFILLER_26_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10810_ _15592_/Q _15591_/Q _15590_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _15584_/D
+ sky130_fd_sc_hd__o31a_1
X_11790_ _11804_/C vssd1 vssd1 vccd1 vccd1 _11814_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ _15574_/Q _10798_/B _10741_/C vssd1 vssd1 vccd1 vccd1 _10750_/B sky130_fd_sc_hd__and3_1
XFILLER_41_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13460_ _13662_/A _13460_/B _13460_/C vssd1 vssd1 vccd1 vccd1 _13462_/B sky130_fd_sc_hd__or3_1
X_10672_ _15563_/Q _10679_/C _10610_/X vssd1 vssd1 vccd1 vccd1 _10672_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ _12636_/A _12414_/C vssd1 vssd1 vccd1 vccd1 _12411_/X sky130_fd_sc_hd__or2_1
X_13391_ _13389_/Y _13384_/C _13387_/X _13388_/Y vssd1 vssd1 vccd1 vccd1 _13392_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _16124_/CLK sky130_fd_sc_hd__clkbuf_16
X_15130_ _15175_/A _15130_/B _15134_/A vssd1 vssd1 vccd1 vccd1 _16351_/D sky130_fd_sc_hd__nor3_1
XFILLER_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ _12350_/A _12340_/Y _12341_/Y _12337_/C vssd1 vssd1 vccd1 vccd1 _12344_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15061_ hold21/X _15131_/B _15061_/C vssd1 vssd1 vccd1 vccd1 _15064_/B sky130_fd_sc_hd__nand3_1
XFILLER_126_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12273_ _12281_/A _12273_/B _12273_/C vssd1 vssd1 vccd1 vccd1 _12274_/A sky130_fd_sc_hd__and3_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14012_ _13912_/X _14010_/B _14011_/Y vssd1 vssd1 vccd1 vccd1 _16104_/D sky130_fd_sc_hd__o21a_1
X_11224_ _11225_/B _11225_/C _11225_/A vssd1 vssd1 vccd1 vccd1 _11226_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11155_ _15646_/Q _15645_/Q _15644_/Q _10983_/X vssd1 vssd1 vccd1 vccd1 _15638_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_122_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10106_ _15475_/Q _10220_/B _10106_/C vssd1 vssd1 vccd1 vccd1 _10115_/B sky130_fd_sc_hd__and3_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11086_ _15628_/Q _11143_/B _11086_/C vssd1 vssd1 vccd1 vccd1 _11094_/B sky130_fd_sc_hd__and3_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15963_ _15984_/CLK _15963_/D vssd1 vssd1 vccd1 vccd1 _15963_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_87_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15259_/CLK sky130_fd_sc_hd__clkbuf_16
X_10037_ _15465_/Q _10155_/B _10037_/C vssd1 vssd1 vccd1 vccd1 _10047_/A sky130_fd_sc_hd__and3_1
X_14914_ _14908_/B _14909_/C _14920_/A _14912_/Y vssd1 vssd1 vccd1 vccd1 _14920_/B
+ sky130_fd_sc_hd__a211oi_1
X_15894_ _07603_/A _15894_/D vssd1 vssd1 vccd1 vccd1 _15894_/Q sky130_fd_sc_hd__dfxtp_1
X_14845_ _15043_/A vssd1 vssd1 vccd1 vccd1 _14845_/X sky130_fd_sc_hd__buf_2
XFILLER_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14776_ _14782_/C vssd1 vssd1 vccd1 vccd1 _14795_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11988_ _11986_/Y _11982_/C _11984_/X _11985_/Y vssd1 vssd1 vccd1 vccd1 _11989_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13727_ _13752_/C vssd1 vssd1 vccd1 vccd1 _13758_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10939_ _15606_/Q _10939_/B _10939_/C vssd1 vssd1 vccd1 vccd1 _10939_/X sky130_fd_sc_hd__and3_1
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13658_ _13658_/A _13658_/B vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12609_/A vssd1 vssd1 vccd1 vccd1 _12840_/B sky130_fd_sc_hd__buf_2
X_13589_ _16032_/Q _13589_/B _13597_/C vssd1 vssd1 vccd1 vccd1 _13589_/X sky130_fd_sc_hd__and3_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _15994_/CLK sky130_fd_sc_hd__clkbuf_16
X_15328_ _15337_/CLK _15328_/D vssd1 vssd1 vccd1 vccd1 _15328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15259_ _15259_/CLK _15259_/D vssd1 vssd1 vccd1 vccd1 _15259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09820_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__nor2_1
X_09751_ _09758_/A _09749_/Y _09750_/Y _09746_/C vssd1 vssd1 vccd1 vccd1 _09753_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15356_/CLK sky130_fd_sc_hd__clkbuf_16
X_08702_ _08699_/X _08700_/Y _08701_/Y _08697_/C vssd1 vssd1 vccd1 vccd1 _08704_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _09680_/Y _09675_/C _09677_/X _09678_/Y vssd1 vssd1 vccd1 vccd1 _09683_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_104_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08633_ _10947_/A vssd1 vssd1 vccd1 vccd1 _13057_/B sky130_fd_sc_hd__buf_4
XFILLER_67_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _08580_/A _08564_/B _08564_/C vssd1 vssd1 vccd1 vccd1 _08565_/A sky130_fd_sc_hd__and3_1
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08495_ _08493_/X _08494_/Y _08488_/B _08489_/C vssd1 vssd1 vccd1 vccd1 _08497_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09116_ _09116_/A vssd1 vssd1 vccd1 vccd1 _15320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09047_ _15310_/Q _09047_/B _09047_/C vssd1 vssd1 vccd1 vccd1 _09047_/Y sky130_fd_sc_hd__nand3_1
XFILLER_108_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09949_ _15451_/Q _09989_/C _09893_/X vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__a21oi_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_69_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15359_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12960_ _12960_/A vssd1 vssd1 vccd1 vccd1 _15922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11911_ _13316_/A vssd1 vssd1 vccd1 vccd1 _13041_/A sky130_fd_sc_hd__buf_2
XFILLER_18_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12906_/A _12891_/B _12891_/C vssd1 vssd1 vccd1 vccd1 _12892_/A sky130_fd_sc_hd__and3_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14630_/A _14630_/B _14630_/C vssd1 vssd1 vccd1 vccd1 _14631_/C sky130_fd_sc_hd__nand3_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11842_/A vssd1 vssd1 vccd1 vccd1 _11883_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14561_/A _14561_/B vssd1 vssd1 vccd1 vccd1 _14561_/Y sky130_fd_sc_hd__nor2_1
X_11773_ _12629_/A vssd1 vssd1 vccd1 vccd1 _12007_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16312_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _16300_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _13662_/A _13512_/B _13512_/C vssd1 vssd1 vccd1 vccd1 _13514_/B sky130_fd_sc_hd__or3_1
X_10724_ _10722_/Y _10718_/C _10720_/X _10721_/Y vssd1 vssd1 vccd1 vccd1 _10725_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14532_/A _14492_/B vssd1 vssd1 vccd1 vccd1 _14493_/B sky130_fd_sc_hd__and2_1
XFILLER_14_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16231_ _16367_/CLK _16231_/D vssd1 vssd1 vccd1 vccd1 _16231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13443_ _13443_/A vssd1 vssd1 vccd1 vccd1 _16003_/D sky130_fd_sc_hd__clkbuf_1
X_10655_ _10940_/A vssd1 vssd1 vccd1 vccd1 _10655_/X sky130_fd_sc_hd__buf_2
XFILLER_139_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16162_ _16166_/CLK _16162_/D vssd1 vssd1 vccd1 vccd1 _16162_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13374_ _15994_/Q _13374_/B _13380_/C vssd1 vssd1 vccd1 vccd1 _13377_/B sky130_fd_sc_hd__nand3_1
X_10586_ _15550_/Q _10623_/C _10474_/X vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__a21oi_1
XFILLER_139_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15113_ _15111_/A _15111_/B _15112_/X vssd1 vssd1 vccd1 vccd1 _16345_/D sky130_fd_sc_hd__a21oi_1
X_12325_ _12609_/A vssd1 vssd1 vccd1 vccd1 _12554_/B sky130_fd_sc_hd__buf_2
XFILLER_115_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16093_ _16103_/CLK _16093_/D vssd1 vssd1 vccd1 vccd1 _16093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15044_ _15038_/A _15041_/B _15043_/X vssd1 vssd1 vccd1 vccd1 _15051_/C sky130_fd_sc_hd__o21a_1
XFILLER_108_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12256_ _15812_/Q _12369_/B _12262_/C vssd1 vssd1 vccd1 vccd1 _12259_/B sky130_fd_sc_hd__nand3_1
X_11207_ _11783_/A vssd1 vssd1 vccd1 vccd1 _11439_/A sky130_fd_sc_hd__clkbuf_2
X_12187_ _12299_/A _12187_/B _12187_/C vssd1 vssd1 vccd1 vccd1 _12190_/B sky130_fd_sc_hd__or3_1
XFILLER_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11138_ _15636_/Q _11143_/C _11137_/X vssd1 vssd1 vccd1 vccd1 _11138_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11069_ _11076_/A _11069_/B _11069_/C vssd1 vssd1 vccd1 vccd1 _11070_/A sky130_fd_sc_hd__and3_1
X_15946_ _15956_/CLK _15946_/D vssd1 vssd1 vccd1 vccd1 _15946_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_0_clk _15665_/CLK vssd1 vssd1 vccd1 vccd1 _15746_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15877_ _15907_/CLK _15877_/D vssd1 vssd1 vccd1 vccd1 _15877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14828_ _14829_/B _14829_/C _14829_/A vssd1 vssd1 vccd1 vccd1 _14830_/B sky130_fd_sc_hd__a21o_1
XFILLER_91_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14759_ _14759_/A _14759_/B vssd1 vssd1 vccd1 vccd1 _14760_/B sky130_fd_sc_hd__nor2_1
X_08280_ _15210_/Q _08403_/B vssd1 vssd1 vccd1 vccd1 _08373_/A sky130_fd_sc_hd__and2_1
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09803_ _15428_/Q _09811_/C _09741_/X vssd1 vssd1 vccd1 vccd1 _09803_/Y sky130_fd_sc_hd__a21oi_1
X_07995_ _16143_/Q vssd1 vssd1 vccd1 vccd1 _14247_/C sky130_fd_sc_hd__inv_2
XFILLER_87_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09734_ _15418_/Q _09735_/C _09506_/X vssd1 vssd1 vccd1 vccd1 _09734_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09665_ _15407_/Q _09721_/B _09671_/C vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__nand3_1
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08616_ _09778_/A vssd1 vssd1 vccd1 vccd1 _08616_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09596_ _10751_/A vssd1 vssd1 vccd1 vccd1 _09596_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _08560_/C vssd1 vssd1 vccd1 vccd1 _08568_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08478_ hold3/X _08532_/C _07623_/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__a21oi_1
XFILLER_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10440_ _15527_/Q _10446_/C _10318_/X vssd1 vssd1 vccd1 vccd1 _10440_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _11582_/A vssd1 vssd1 vccd1 vccd1 _10602_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_124_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _12107_/X _12108_/Y _12109_/Y _12105_/C vssd1 vssd1 vccd1 vccd1 _12112_/B
+ sky130_fd_sc_hd__o211ai_1
X_13090_ _15962_/Q _15961_/Q _15960_/Q _12981_/X vssd1 vssd1 vccd1 vccd1 _15945_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_105_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12041_ _12041_/A vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15800_ _15809_/CLK _15800_/D vssd1 vssd1 vccd1 vccd1 _15800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13992_ _13998_/A _13991_/Y _13985_/B _13986_/C vssd1 vssd1 vccd1 vccd1 _13994_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15731_ _15794_/CLK _15731_/D vssd1 vssd1 vccd1 vccd1 _15731_/Q sky130_fd_sc_hd__dfxtp_1
X_12943_ _12941_/X _12942_/Y _12938_/B _12939_/C vssd1 vssd1 vccd1 vccd1 _12945_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15662_ _15763_/CLK _15662_/D vssd1 vssd1 vccd1 vccd1 _15662_/Q sky130_fd_sc_hd__dfxtp_1
X_12874_ _12874_/A vssd1 vssd1 vccd1 vccd1 _12887_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _11825_/A vssd1 vssd1 vccd1 vccd1 _15742_/D sky130_fd_sc_hd__clkbuf_1
X_14613_ _07688_/X _14611_/B _14612_/Y vssd1 vssd1 vccd1 vccd1 _16230_/D sky130_fd_sc_hd__o21a_1
X_15593_ _15602_/CLK _15593_/D vssd1 vssd1 vccd1 vccd1 _15593_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14554_/C vssd1 vssd1 vccd1 vccd1 _14566_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11756_ _11754_/Y _11749_/C _11751_/X _11752_/Y vssd1 vssd1 vccd1 vccd1 _11757_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10707_ _15569_/Q _10876_/B _10714_/C vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__nand3_1
XFILLER_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14475_ _16203_/Q _14474_/C _14300_/X vssd1 vssd1 vccd1 vccd1 _14475_/Y sky130_fd_sc_hd__a21oi_1
X_11687_ _11708_/A _11687_/B _11687_/C vssd1 vssd1 vccd1 vccd1 _11688_/A sky130_fd_sc_hd__and3_1
X_13426_ _13427_/B _13427_/C _13427_/A vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__a21o_1
X_16214_ _16222_/CLK _16214_/D vssd1 vssd1 vccd1 vccd1 _16214_/Q sky130_fd_sc_hd__dfxtp_1
X_10638_ _15565_/Q _15564_/Q _15563_/Q _10409_/X vssd1 vssd1 vccd1 vccd1 _15557_/D
+ sky130_fd_sc_hd__o31a_1
X_16145_ _16148_/CLK _16145_/D vssd1 vssd1 vccd1 vccd1 _16145_/Q sky130_fd_sc_hd__dfxtp_2
X_13357_ _13612_/A vssd1 vssd1 vccd1 vccd1 _13410_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10569_ _15547_/Q _10798_/B _10569_/C vssd1 vssd1 vccd1 vccd1 _10577_/B sky130_fd_sc_hd__and3_1
XFILLER_127_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12308_ _15820_/Q _12346_/C _12197_/X vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__a21oi_1
XFILLER_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16076_ _16143_/CLK _16076_/D vssd1 vssd1 vccd1 vccd1 _16076_/Q sky130_fd_sc_hd__dfxtp_1
X_13288_ _13286_/Y _13281_/C _13284_/X _13285_/Y vssd1 vssd1 vccd1 vccd1 _13289_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_114_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15027_ _15027_/A _15027_/B _15027_/C vssd1 vssd1 vccd1 vccd1 _15028_/C sky130_fd_sc_hd__nand3_1
X_12239_ _12239_/A _12239_/B vssd1 vssd1 vccd1 vccd1 _12243_/C sky130_fd_sc_hd__nor2_1
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07780_ _07780_/A _07780_/B vssd1 vssd1 vccd1 vccd1 _07781_/B sky130_fd_sc_hd__xor2_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 in1[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_8
XFILLER_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15929_ _15196_/Q _15929_/D vssd1 vssd1 vccd1 vccd1 _15929_/Q sky130_fd_sc_hd__dfxtp_1
X_09450_ _09450_/A vssd1 vssd1 vccd1 vccd1 _15372_/D sky130_fd_sc_hd__clkbuf_1
X_08401_ _08401_/A vssd1 vssd1 vccd1 vccd1 _15211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09381_ _15363_/Q _09391_/C _09212_/X vssd1 vssd1 vccd1 vccd1 _09381_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08332_ _08436_/A _08332_/B vssd1 vssd1 vccd1 vccd1 _08332_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08263_ _08263_/A _08263_/B vssd1 vssd1 vccd1 vccd1 _08266_/A sky130_fd_sc_hd__xnor2_4
XFILLER_137_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08194_ _08194_/A _08292_/A vssd1 vssd1 vccd1 vccd1 _08287_/A sky130_fd_sc_hd__xor2_4
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07978_ _08195_/B _07978_/B vssd1 vssd1 vccd1 vccd1 _07979_/B sky130_fd_sc_hd__xnor2_2
X_09717_ _15415_/Q _09754_/C _09605_/X vssd1 vssd1 vccd1 vccd1 _09720_/B sky130_fd_sc_hd__a21oi_1
XFILLER_68_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09648_ _09648_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09652_/C sky130_fd_sc_hd__nor2_1
XFILLER_55_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _11080_/A vssd1 vssd1 vccd1 vccd1 _10736_/A sky130_fd_sc_hd__buf_2
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11780_/A _11614_/C vssd1 vssd1 vccd1 vccd1 _11610_/X sky130_fd_sc_hd__or2_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12590_ _12610_/C vssd1 vssd1 vccd1 vccd1 _12623_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11541_ _15699_/Q _11655_/B _11541_/C vssd1 vssd1 vccd1 vccd1 _11550_/A sky130_fd_sc_hd__and3_1
XFILLER_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14260_ _14304_/A _14260_/B _14264_/B vssd1 vssd1 vccd1 vccd1 _16155_/D sky130_fd_sc_hd__nor3_1
XFILLER_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _12048_/A vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13211_ _15954_/Q vssd1 vssd1 vccd1 vccd1 _13217_/C sky130_fd_sc_hd__inv_2
X_10423_ _10423_/A vssd1 vssd1 vccd1 vccd1 _15523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14191_ _14183_/Y _14185_/X _14187_/B vssd1 vssd1 vccd1 vccd1 _14192_/B sky130_fd_sc_hd__o21a_1
XFILLER_124_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13142_ _13142_/A _13142_/B vssd1 vssd1 vccd1 vccd1 _13146_/C sky130_fd_sc_hd__nor2_1
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10354_ _10354_/A vssd1 vssd1 vccd1 vccd1 _11569_/A sky130_fd_sc_hd__buf_4
XFILLER_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13073_ _13700_/A vssd1 vssd1 vccd1 vccd1 _14402_/A sky130_fd_sc_hd__clkbuf_4
X_10285_ _10284_/B _10284_/C _10172_/X vssd1 vssd1 vccd1 vccd1 _10286_/C sky130_fd_sc_hd__o21ai_1
X_12024_ _15775_/Q _12062_/C _11912_/X vssd1 vssd1 vccd1 vccd1 _12026_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13975_ _16089_/Q vssd1 vssd1 vccd1 vccd1 _13979_/C sky130_fd_sc_hd__inv_2
XFILLER_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15714_ _15794_/CLK _15714_/D vssd1 vssd1 vccd1 vccd1 _15714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _12926_/A vssd1 vssd1 vccd1 vccd1 _15916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15645_ _15655_/CLK _15645_/D vssd1 vssd1 vccd1 vccd1 _15645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _15905_/Q _13018_/B _12861_/C vssd1 vssd1 vccd1 vccd1 _12857_/Y sky130_fd_sc_hd__nand3_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _11801_/B _11802_/C _11804_/X _11806_/Y vssd1 vssd1 vccd1 vccd1 _11809_/C
+ sky130_fd_sc_hd__a211o_1
X_15576_ _15194_/Q _15576_/D vssd1 vssd1 vccd1 vccd1 _15576_/Q sky130_fd_sc_hd__dfxtp_2
X_12788_ _12786_/Y _12782_/C _12784_/X _12785_/Y vssd1 vssd1 vccd1 vccd1 _12789_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11739_ _15731_/Q _11797_/B _11745_/C vssd1 vssd1 vccd1 vccd1 _11742_/B sky130_fd_sc_hd__nand3_1
X_14527_ _14525_/X _14527_/B vssd1 vssd1 vccd1 vccd1 _14527_/X sky130_fd_sc_hd__and2b_1
XFILLER_30_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14458_ _14325_/X _14454_/B _14326_/X vssd1 vssd1 vccd1 vccd1 _14461_/A sky130_fd_sc_hd__a21oi_1
XFILLER_127_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13409_ _13408_/B _13408_/C _13305_/X vssd1 vssd1 vccd1 vccd1 _13410_/C sky130_fd_sc_hd__o21ai_1
X_14389_ _16185_/Q _14474_/B _14389_/C vssd1 vssd1 vccd1 vccd1 _14397_/A sky130_fd_sc_hd__and3_1
XFILLER_142_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16128_ _16129_/CLK _16128_/D vssd1 vssd1 vccd1 vccd1 _16128_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08950_ _09066_/A _08950_/B _08954_/B vssd1 vssd1 vccd1 vccd1 _15294_/D sky130_fd_sc_hd__nor3_1
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16059_ _16075_/CLK _16059_/D vssd1 vssd1 vccd1 vccd1 _16059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07901_ _16179_/Q _16197_/Q vssd1 vssd1 vccd1 vccd1 _07967_/B sky130_fd_sc_hd__xor2_4
X_08881_ _15286_/Q _08886_/C _08824_/X vssd1 vssd1 vccd1 vccd1 _08881_/Y sky130_fd_sc_hd__a21oi_1
X_07832_ _15638_/Q vssd1 vssd1 vccd1 vccd1 _11156_/A sky130_fd_sc_hd__clkinv_2
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07763_ _15503_/Q _15485_/Q vssd1 vssd1 vccd1 vccd1 _08093_/B sky130_fd_sc_hd__xor2_4
X_09502_ _09502_/A vssd1 vssd1 vccd1 vccd1 _15380_/D sky130_fd_sc_hd__clkbuf_1
X_07694_ _10969_/A vssd1 vssd1 vccd1 vccd1 _12631_/A sky130_fd_sc_hd__clkbuf_4
X_09433_ _15371_/Q _09438_/C _09205_/X vssd1 vssd1 vccd1 vccd1 _09435_/C sky130_fd_sc_hd__a21o_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09401_/A _09364_/B _09364_/C vssd1 vssd1 vccd1 vccd1 _09365_/A sky130_fd_sc_hd__and3_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08315_ _08315_/A _08315_/B vssd1 vssd1 vccd1 vccd1 _08316_/B sky130_fd_sc_hd__nand2_1
XANTENNA_20 _13720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09295_ _09293_/Y _09288_/C _09300_/A _09291_/Y vssd1 vssd1 vccd1 vccd1 _09300_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA_31 _14988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08246_ _08246_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _08246_/X sky130_fd_sc_hd__or2_1
XFILLER_119_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08177_ _08177_/A _07984_/A vssd1 vssd1 vccd1 vccd1 _08179_/A sky130_fd_sc_hd__or2b_1
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10070_ _10071_/B _10071_/C _10071_/A vssd1 vssd1 vccd1 vccd1 _10072_/B sky130_fd_sc_hd__a21o_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ _13766_/B _13760_/B vssd1 vssd1 vccd1 vccd1 _13763_/A sky130_fd_sc_hd__or2_1
X_10972_ _10979_/B _10972_/B vssd1 vssd1 vccd1 vccd1 _10975_/A sky130_fd_sc_hd__or2_1
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ _15883_/Q _12879_/B _12720_/C vssd1 vssd1 vccd1 vccd1 _12717_/A sky130_fd_sc_hd__and3_1
X_13691_ _13691_/A vssd1 vssd1 vccd1 vccd1 _16047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15430_ _15484_/CLK _15430_/D vssd1 vssd1 vccd1 vccd1 _15430_/Q sky130_fd_sc_hd__dfxtp_1
X_12642_ _12680_/A _12642_/B _12642_/C vssd1 vssd1 vccd1 vccd1 _12643_/A sky130_fd_sc_hd__and3_1
XFILLER_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15361_ _15377_/CLK _15361_/D vssd1 vssd1 vccd1 vccd1 _15361_/Q sky130_fd_sc_hd__dfxtp_1
X_12573_ _12571_/Y _12565_/C _12578_/A _12570_/Y vssd1 vssd1 vccd1 vccd1 _12578_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14312_ _14308_/B _14307_/Y _14308_/A vssd1 vssd1 vccd1 vccd1 _14312_/Y sky130_fd_sc_hd__o21bai_1
X_11524_ _11524_/A vssd1 vssd1 vccd1 vccd1 _15695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15292_ _15301_/CLK _15292_/D vssd1 vssd1 vccd1 vccd1 _15292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14243_ _16169_/Q _16168_/Q _16167_/Q _14202_/X vssd1 vssd1 vccd1 vccd1 _16152_/D
+ sky130_fd_sc_hd__o31a_1
X_11455_ _11477_/A _11455_/B _11455_/C vssd1 vssd1 vccd1 vccd1 _11456_/A sky130_fd_sc_hd__and3_1
XFILLER_125_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10406_ _10405_/B _10405_/C _10172_/X vssd1 vssd1 vccd1 vccd1 _10407_/C sky130_fd_sc_hd__o21ai_1
XFILLER_124_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14174_ _14168_/B _14169_/C _14179_/A _14172_/Y vssd1 vssd1 vccd1 vccd1 _14179_/B
+ sky130_fd_sc_hd__a211oi_1
X_11386_ _15682_/Q _15681_/Q _15680_/Q _11273_/X vssd1 vssd1 vccd1 vccd1 _15674_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_98_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ _13149_/A _13125_/B _13125_/C vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__and3_1
X_10337_ _10337_/A _10337_/B vssd1 vssd1 vccd1 vccd1 _10342_/C sky130_fd_sc_hd__nor2_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13056_/A vssd1 vssd1 vccd1 vccd1 _15939_/D sky130_fd_sc_hd__clkbuf_1
X_10268_ _15501_/Q _10446_/B _10268_/C vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__and3_1
XFILLER_140_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12007_ _15772_/Q _12007_/B _12007_/C vssd1 vssd1 vccd1 vccd1 _12015_/B sky130_fd_sc_hd__and3_1
X_10199_ _15489_/Q _10199_/B _10199_/C vssd1 vssd1 vccd1 vccd1 _10199_/Y sky130_fd_sc_hd__nand3_1
XFILLER_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13958_ _16097_/Q _13957_/C _15043_/A vssd1 vssd1 vccd1 vccd1 _13959_/B sky130_fd_sc_hd__a21o_1
X_12909_ _15915_/Q _12914_/C _12855_/X vssd1 vssd1 vccd1 vccd1 _12909_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13889_ _13980_/A _13889_/B _13895_/B vssd1 vssd1 vccd1 vccd1 _16083_/D sky130_fd_sc_hd__nor3_1
XFILLER_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15628_ _15194_/Q _15628_/D vssd1 vssd1 vccd1 vccd1 _15628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ _15655_/CLK _15559_/D vssd1 vssd1 vccd1 vccd1 _15559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08100_ _14863_/C _08100_/B vssd1 vssd1 vccd1 vccd1 _08100_/X sky130_fd_sc_hd__or2_1
X_09080_ _13930_/A vssd1 vssd1 vccd1 vccd1 _11963_/A sky130_fd_sc_hd__buf_6
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08031_ _12588_/A _12706_/A _08030_/Y vssd1 vssd1 vccd1 vccd1 _08033_/C sky130_fd_sc_hd__o21a_1
XFILLER_135_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09982_ _15456_/Q _09989_/C _09981_/X vssd1 vssd1 vccd1 vccd1 _09982_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08933_ _08931_/Y _08924_/C _08928_/X _08930_/Y vssd1 vssd1 vccd1 vccd1 _08934_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08864_ _08864_/A vssd1 vssd1 vccd1 vccd1 _15282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07815_ _15791_/Q _08052_/A _07815_/C vssd1 vssd1 vccd1 vccd1 _08052_/B sky130_fd_sc_hd__nand3_1
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08795_ _08909_/A _08795_/B _08799_/A vssd1 vssd1 vccd1 vccd1 _15271_/D sky130_fd_sc_hd__nor3_1
XFILLER_123_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07746_ _08106_/A _08107_/B vssd1 vssd1 vccd1 vccd1 _07752_/A sky130_fd_sc_hd__xnor2_4
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07677_ _07665_/A _07668_/B _15001_/A vssd1 vssd1 vccd1 vccd1 _07698_/C sky130_fd_sc_hd__o21a_1
XFILLER_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09416_ _09472_/A _09419_/C vssd1 vssd1 vccd1 vccd1 _09416_/X sky130_fd_sc_hd__or2_1
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09347_ _09924_/A vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__buf_2
XFILLER_32_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ _15346_/Q _09334_/B _09278_/C vssd1 vssd1 vccd1 vccd1 _09278_/Y sky130_fd_sc_hd__nand3_1
XFILLER_138_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ _08075_/A _08075_/B _08228_/Y vssd1 vssd1 vccd1 vccd1 _08231_/C sky130_fd_sc_hd__a21oi_1
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _11236_/X _11238_/Y _11239_/Y _11234_/C vssd1 vssd1 vccd1 vccd1 _11242_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_146_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11171_ _11169_/X _11170_/Y _11166_/B _11167_/C vssd1 vssd1 vccd1 vccd1 _11173_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10122_ _10135_/C vssd1 vssd1 vccd1 vccd1 _10143_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10053_ _10284_/A _10053_/B _10053_/C vssd1 vssd1 vccd1 vccd1 _10055_/B sky130_fd_sc_hd__or3_1
X_14930_ _15051_/A _15010_/B _14930_/C vssd1 vssd1 vccd1 vccd1 _14932_/A sky130_fd_sc_hd__and3_1
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14861_ _16292_/Q _14977_/B _14863_/C vssd1 vssd1 vccd1 vccd1 _14866_/A sky130_fd_sc_hd__and3_1
XFILLER_91_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13812_ _14106_/A _13812_/B _13812_/C vssd1 vssd1 vccd1 vccd1 _13814_/B sky130_fd_sc_hd__or3_1
XFILLER_90_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14792_ _14785_/B _14786_/C _14798_/A _14790_/Y vssd1 vssd1 vccd1 vccd1 _14798_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13743_ _13743_/A vssd1 vssd1 vccd1 vccd1 _16056_/D sky130_fd_sc_hd__clkbuf_1
X_10955_ _15608_/Q _10963_/B _11080_/A vssd1 vssd1 vccd1 vccd1 _10955_/X sky130_fd_sc_hd__and3_1
XFILLER_44_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13674_ _16047_/Q _13707_/C _13573_/X vssd1 vssd1 vccd1 vccd1 _13676_/B sky130_fd_sc_hd__a21oi_1
X_10886_ _10902_/A _10886_/B _10886_/C vssd1 vssd1 vccd1 vccd1 _10887_/A sky130_fd_sc_hd__and3_1
XFILLER_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15413_ _15422_/CLK _15413_/D vssd1 vssd1 vccd1 vccd1 _15413_/Q sky130_fd_sc_hd__dfxtp_2
X_12625_ _15869_/Q _12744_/B _12630_/C vssd1 vssd1 vccd1 vccd1 _12625_/Y sky130_fd_sc_hd__nand3_1
X_15344_ _15348_/CLK _15344_/D vssd1 vssd1 vccd1 vccd1 _15344_/Q sky130_fd_sc_hd__dfxtp_1
X_12556_ _12554_/Y _12550_/C _12552_/X _12553_/Y vssd1 vssd1 vccd1 vccd1 _12557_/C
+ sky130_fd_sc_hd__a211o_1
X_11507_ _11507_/A vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15275_ _15286_/CLK _15275_/D vssd1 vssd1 vccd1 vccd1 _15275_/Q sky130_fd_sc_hd__dfxtp_1
X_12487_ _12488_/B _12488_/C _12488_/A vssd1 vssd1 vccd1 vccd1 _12489_/B sky130_fd_sc_hd__a21o_1
XFILLER_144_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14226_ _14224_/A _14224_/B _14223_/Y _14225_/Y vssd1 vssd1 vccd1 vccd1 _16147_/D
+ sky130_fd_sc_hd__o31a_1
X_11438_ _11555_/A vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14157_ _14161_/C vssd1 vssd1 vccd1 vccd1 _14171_/C sky130_fd_sc_hd__clkbuf_1
X_11369_ _12230_/A vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_140_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13108_ _13532_/A vssd1 vssd1 vccd1 vccd1 _14298_/A sky130_fd_sc_hd__buf_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _16121_/Q _14088_/B _14093_/C vssd1 vssd1 vccd1 vccd1 _14088_/Y sky130_fd_sc_hd__nand3_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _13059_/C vssd1 vssd1 vccd1 vccd1 _13071_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07600_ _08944_/A vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__buf_4
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08580_ _08580_/A _08580_/B _08580_/C vssd1 vssd1 vccd1 vccd1 _08581_/A sky130_fd_sc_hd__and3_1
XFILLER_93_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09201_ _15335_/Q _09372_/B _09211_/C vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__and3_1
XFILLER_50_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09132_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09171_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ _15312_/Q _09238_/B _09067_/C vssd1 vssd1 vccd1 vccd1 _09063_/Y sky130_fd_sc_hd__nand3_1
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08014_ _08014_/A _08014_/B vssd1 vssd1 vccd1 vccd1 _08205_/B sky130_fd_sc_hd__xnor2_1
XFILLER_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09965_ _15454_/Q _09967_/C _09794_/X vssd1 vssd1 vccd1 vccd1 _09965_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08916_ _08916_/A _08916_/B _08916_/C vssd1 vssd1 vccd1 vccd1 _08917_/C sky130_fd_sc_hd__nand3_1
X_09896_ _09930_/A _09896_/B _09900_/A vssd1 vssd1 vccd1 vccd1 _15441_/D sky130_fd_sc_hd__nor3_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08847_ _08880_/C vssd1 vssd1 vccd1 vccd1 _08886_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08778_ _08778_/A _08778_/B vssd1 vssd1 vccd1 vccd1 _08779_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07729_ _07729_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _08132_/B sky130_fd_sc_hd__xor2_4
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ _10797_/A _10740_/B _10744_/B vssd1 vssd1 vccd1 vccd1 _15572_/D sky130_fd_sc_hd__nor3_1
XFILLER_81_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10671_ _15563_/Q _10895_/B _10679_/C vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__and3_1
XFILLER_41_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12410_ _12410_/A _12410_/B vssd1 vssd1 vccd1 vccd1 _12414_/C sky130_fd_sc_hd__nor2_1
X_13390_ _13387_/X _13388_/Y _13389_/Y _13384_/C vssd1 vssd1 vccd1 vccd1 _13392_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12341_ _15824_/Q _12458_/B _12346_/C vssd1 vssd1 vccd1 vccd1 _12341_/Y sky130_fd_sc_hd__nand3_1
XFILLER_139_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15060_ _15106_/A _15060_/B _15064_/A vssd1 vssd1 vccd1 vccd1 _16333_/D sky130_fd_sc_hd__nor3_1
X_12272_ _12270_/Y _12266_/C _12268_/X _12269_/Y vssd1 vssd1 vccd1 vccd1 _12273_/C
+ sky130_fd_sc_hd__a211o_1
X_14011_ _14054_/A _14011_/B vssd1 vssd1 vccd1 vccd1 _14011_/Y sky130_fd_sc_hd__nor2_1
X_11223_ _15650_/Q _11228_/C _11222_/X vssd1 vssd1 vccd1 vccd1 _11225_/C sky130_fd_sc_hd__a21o_1
XFILLER_135_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11154_ _11154_/A vssd1 vssd1 vccd1 vccd1 _15637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10105_ _10219_/A _10105_/B _10109_/B vssd1 vssd1 vccd1 vccd1 _15473_/D sky130_fd_sc_hd__nor3_1
X_11085_ _11085_/A _11085_/B _11089_/B vssd1 vssd1 vccd1 vccd1 _15626_/D sky130_fd_sc_hd__nor3_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15962_ _15971_/CLK _15962_/D vssd1 vssd1 vccd1 vccd1 _15962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10036_ _10036_/A vssd1 vssd1 vccd1 vccd1 _15463_/D sky130_fd_sc_hd__clkbuf_1
X_14913_ _14920_/A _14912_/Y _14908_/B _14909_/C vssd1 vssd1 vccd1 vccd1 _14915_/B
+ sky130_fd_sc_hd__o211a_1
X_15893_ _07603_/A _15893_/D vssd1 vssd1 vccd1 vccd1 _15893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14844_ _14842_/A _14842_/B _14843_/X vssd1 vssd1 vccd1 vccd1 _16282_/D sky130_fd_sc_hd__a21oi_1
XFILLER_17_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14775_ _16286_/Q _16285_/Q _16284_/Q _14620_/X vssd1 vssd1 vccd1 vccd1 _16269_/D
+ sky130_fd_sc_hd__o31a_1
X_11987_ _11984_/X _11985_/Y _11986_/Y _11982_/C vssd1 vssd1 vccd1 vccd1 _11989_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13726_ _13738_/C vssd1 vssd1 vccd1 vccd1 _13752_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10938_ _10938_/A vssd1 vssd1 vccd1 vccd1 _15604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10869_ _10882_/C vssd1 vssd1 vccd1 vccd1 _10890_/C sky130_fd_sc_hd__clkbuf_1
X_13657_ _13662_/B _13657_/B vssd1 vssd1 vccd1 vccd1 _13659_/A sky130_fd_sc_hd__or2_1
XFILLER_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12608_ _15868_/Q _12610_/C _12384_/X vssd1 vssd1 vccd1 vccd1 _12608_/Y sky130_fd_sc_hd__a21oi_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13588_ _13588_/A vssd1 vssd1 vccd1 vccd1 _16029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15327_ _15337_/CLK _15327_/D vssd1 vssd1 vccd1 vccd1 _15327_/Q sky130_fd_sc_hd__dfxtp_1
X_12539_ _12652_/A _12539_/B _12543_/A vssd1 vssd1 vccd1 vccd1 _15855_/D sky130_fd_sc_hd__nor3_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15258_ _15259_/CLK _15258_/D vssd1 vssd1 vccd1 vccd1 _15258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14209_ _16148_/Q _14249_/B _14216_/C vssd1 vssd1 vccd1 vccd1 _14212_/B sky130_fd_sc_hd__nand3_1
XFILLER_125_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15189_ _15189_/A _15189_/B _15189_/C vssd1 vssd1 vccd1 vccd1 _15191_/A sky130_fd_sc_hd__and3_1
XFILLER_125_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09750_ _15419_/Q _09813_/B _09754_/C vssd1 vssd1 vccd1 vccd1 _09750_/Y sky130_fd_sc_hd__nand3_1
XFILLER_101_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08701_ _15257_/Q _10957_/C _08706_/C vssd1 vssd1 vccd1 vccd1 _08701_/Y sky130_fd_sc_hd__nand3_1
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09681_ _09677_/X _09678_/Y _09680_/Y _09675_/C vssd1 vssd1 vccd1 vccd1 _09683_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_55_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08632_ _15248_/Q _08865_/B _08636_/C vssd1 vssd1 vccd1 vccd1 _08632_/X sky130_fd_sc_hd__and3_1
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08563_ _08557_/B _08558_/C _08560_/X _08561_/Y vssd1 vssd1 vccd1 vccd1 _08564_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _15229_/Q _08505_/C _12609_/A vssd1 vssd1 vccd1 vccd1 _08494_/Y sky130_fd_sc_hd__a21oi_1
X_09115_ _09115_/A _09115_/B _09115_/C vssd1 vssd1 vccd1 vccd1 _09116_/A sky130_fd_sc_hd__and3_1
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09046_ _15311_/Q _09047_/C _08929_/X vssd1 vssd1 vccd1 vccd1 _09046_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09948_ _09979_/C vssd1 vssd1 vccd1 vccd1 _09989_/C sky130_fd_sc_hd__clkbuf_2
X_09879_ _10049_/A _09883_/C vssd1 vssd1 vccd1 vccd1 _09879_/X sky130_fd_sc_hd__or2_1
XFILLER_46_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11910_ _11943_/C vssd1 vssd1 vccd1 vccd1 _11950_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_100_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12890_ _12884_/B _12885_/C _12887_/X _12888_/Y vssd1 vssd1 vccd1 vccd1 _12891_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11839_/A _11839_/B _11840_/X vssd1 vssd1 vccd1 vccd1 _15744_/D sky130_fd_sc_hd__a21oi_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11796_/A _11772_/B _11778_/B vssd1 vssd1 vccd1 vccd1 _15734_/D sky130_fd_sc_hd__nor3_1
XFILLER_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14560_ _16222_/Q _14566_/C _14395_/X vssd1 vssd1 vccd1 vccd1 _14562_/B sky130_fd_sc_hd__a21oi_1
XFILLER_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _10720_/X _10721_/Y _10722_/Y _10718_/C vssd1 vssd1 vccd1 vccd1 _10725_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13509_/A _13509_/B _13510_/X vssd1 vssd1 vccd1 vccd1 _16014_/D sky130_fd_sc_hd__a21oi_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _14485_/Y _14486_/X _14488_/B vssd1 vssd1 vccd1 vccd1 _14492_/B sky130_fd_sc_hd__o21a_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16230_ _16362_/CLK _16230_/D vssd1 vssd1 vccd1 vccd1 _16230_/Q sky130_fd_sc_hd__dfxtp_1
X_10654_ _15561_/Q _10654_/B _10654_/C vssd1 vssd1 vccd1 vccd1 _10654_/X sky130_fd_sc_hd__and3_1
X_13442_ _13481_/A _13442_/B _13442_/C vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__and3_1
XFILLER_9_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13373_ _13476_/A _13373_/B _13377_/A vssd1 vssd1 vccd1 vccd1 _15991_/D sky130_fd_sc_hd__nor3_1
X_16161_ _16187_/CLK _16161_/D vssd1 vssd1 vccd1 vccd1 _16161_/Q sky130_fd_sc_hd__dfxtp_2
X_10585_ _10617_/C vssd1 vssd1 vccd1 vccd1 _10623_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15112_ _15181_/A _15112_/B vssd1 vssd1 vccd1 vccd1 _15112_/X sky130_fd_sc_hd__or2_1
X_12324_ _15823_/Q _12326_/C _12100_/X vssd1 vssd1 vccd1 vccd1 _12324_/Y sky130_fd_sc_hd__a21oi_1
X_16092_ _16224_/CLK _16092_/D vssd1 vssd1 vccd1 vccd1 _16092_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12255_ _12368_/A _12255_/B _12259_/A vssd1 vssd1 vccd1 vccd1 _15810_/D sky130_fd_sc_hd__nor3_1
X_15043_ _15043_/A vssd1 vssd1 vccd1 vccd1 _15043_/X sky130_fd_sc_hd__buf_2
XFILLER_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11206_ _11267_/A vssd1 vssd1 vccd1 vccd1 _11249_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12186_ _12413_/A vssd1 vssd1 vccd1 vccd1 _12226_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11137_ _11137_/A vssd1 vssd1 vccd1 vccd1 _11137_/X sky130_fd_sc_hd__buf_2
XFILLER_96_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11068_ _11066_/Y _11062_/C _11064_/X _11065_/Y vssd1 vssd1 vccd1 vccd1 _11069_/C
+ sky130_fd_sc_hd__a211o_1
X_15945_ _15970_/CLK _15945_/D vssd1 vssd1 vccd1 vccd1 _15945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10019_ _10013_/B _10014_/C _10016_/X _10017_/Y vssd1 vssd1 vccd1 vccd1 _10020_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_37_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15876_ _07603_/A _15876_/D vssd1 vssd1 vccd1 vccd1 _15876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14827_ _16284_/Q _14826_/C _14744_/X vssd1 vssd1 vccd1 vccd1 _14829_/C sky130_fd_sc_hd__a21o_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16369__18 vssd1 vssd1 vccd1 vccd1 _16369__18/HI io_oeb[1] sky130_fd_sc_hd__conb_1
X_14758_ _14758_/A _14758_/B vssd1 vssd1 vccd1 vccd1 _14759_/B sky130_fd_sc_hd__nor2_1
X_13709_ _16052_/Q _13707_/C _13708_/X vssd1 vssd1 vccd1 vccd1 _13710_/B sky130_fd_sc_hd__a21oi_1
X_14689_ _14765_/A _14693_/C vssd1 vssd1 vccd1 vccd1 _14691_/A sky130_fd_sc_hd__and2_1
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16359_ _16359_/CLK _16359_/D vssd1 vssd1 vccd1 vccd1 _16359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09802_ _15428_/Q _10029_/B _09811_/C vssd1 vssd1 vccd1 vccd1 _09802_/X sky130_fd_sc_hd__and3_1
XFILLER_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07994_ _16125_/Q vssd1 vssd1 vccd1 vccd1 _14161_/C sky130_fd_sc_hd__inv_2
XFILLER_87_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09733_ _15418_/Q _09733_/B _09735_/C vssd1 vssd1 vccd1 vccd1 _09733_/X sky130_fd_sc_hd__and3_1
XFILLER_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09664_ _09775_/A _09664_/B _09668_/A vssd1 vssd1 vccd1 vccd1 _15405_/D sky130_fd_sc_hd__nor3_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08615_ _10354_/A vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__clkbuf_8
X_09595_ _11037_/A vssd1 vssd1 vccd1 vccd1 _10751_/A sky130_fd_sc_hd__buf_4
XFILLER_55_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _08546_/A vssd1 vssd1 vccd1 vccd1 _08560_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08477_ _08522_/C vssd1 vssd1 vccd1 vccd1 _08532_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10370_ input4/X vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__buf_4
XFILLER_108_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09029_ _10181_/A vssd1 vssd1 vccd1 vccd1 _09029_/X sky130_fd_sc_hd__buf_2
XFILLER_108_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _15778_/Q _12042_/C _11812_/X vssd1 vssd1 vccd1 vccd1 _12040_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13991_ _16104_/Q _13990_/C _14088_/B vssd1 vssd1 vccd1 vccd1 _13991_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15730_ _15794_/CLK _15730_/D vssd1 vssd1 vccd1 vccd1 _15730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12942_ _15921_/Q _12949_/C _13275_/A vssd1 vssd1 vccd1 vccd1 _12942_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15661_ _15763_/CLK _15661_/D vssd1 vssd1 vccd1 vccd1 _15661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12873_ _15914_/Q _15916_/Q _15915_/Q _12704_/X vssd1 vssd1 vccd1 vccd1 _15908_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14612_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14612_/Y sky130_fd_sc_hd__nor2_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _11824_/A _11824_/B _11824_/C vssd1 vssd1 vccd1 vccd1 _11825_/A sky130_fd_sc_hd__and3_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15194_/Q _15592_/D vssd1 vssd1 vccd1 vccd1 _15592_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _14546_/C vssd1 vssd1 vccd1 vccd1 _14554_/C sky130_fd_sc_hd__clkbuf_1
X_11755_ _11751_/X _11752_/Y _11754_/Y _11749_/C vssd1 vssd1 vccd1 vccd1 _11757_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_42_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _10797_/A _10706_/B _10710_/A vssd1 vssd1 vccd1 vccd1 _15567_/D sky130_fd_sc_hd__nor3_1
X_14474_ _16203_/Q _14474_/B _14474_/C vssd1 vssd1 vccd1 vccd1 _14481_/A sky130_fd_sc_hd__and3_1
X_11686_ _11686_/A _11686_/B _11686_/C vssd1 vssd1 vccd1 vccd1 _11687_/C sky130_fd_sc_hd__nand3_1
X_16213_ _16222_/CLK _16213_/D vssd1 vssd1 vccd1 vccd1 _16213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13425_ _16003_/Q _13430_/C _13269_/X vssd1 vssd1 vccd1 vccd1 _13427_/C sky130_fd_sc_hd__a21o_1
X_10637_ _10637_/A vssd1 vssd1 vccd1 vccd1 _15556_/D sky130_fd_sc_hd__clkbuf_1
X_16144_ _16148_/CLK _16144_/D vssd1 vssd1 vccd1 vccd1 _16144_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10568_ _11197_/A vssd1 vssd1 vccd1 vccd1 _10798_/B sky130_fd_sc_hd__clkbuf_2
X_13356_ _14163_/A vssd1 vssd1 vccd1 vccd1 _13612_/A sky130_fd_sc_hd__buf_2
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ _12339_/C vssd1 vssd1 vccd1 vccd1 _12346_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_114_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16075_ _16075_/CLK _16075_/D vssd1 vssd1 vccd1 vccd1 _16075_/Q sky130_fd_sc_hd__dfxtp_1
X_10499_ _10785_/A vssd1 vssd1 vccd1 vccd1 _10729_/B sky130_fd_sc_hd__buf_2
XFILLER_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13287_ _13284_/X _13285_/Y _13286_/Y _13281_/C vssd1 vssd1 vccd1 vccd1 _13289_/B
+ sky130_fd_sc_hd__o211ai_1
X_15026_ _15027_/B _15027_/C _15027_/A vssd1 vssd1 vccd1 vccd1 _15028_/B sky130_fd_sc_hd__a21o_1
X_12238_ _12238_/A _12238_/B vssd1 vssd1 vccd1 vccd1 _12239_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _12167_/Y _12162_/C _12165_/X _12166_/Y vssd1 vssd1 vccd1 vccd1 _12170_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 in1[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
X_15928_ _15196_/Q _15928_/D vssd1 vssd1 vccd1 vccd1 _15928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15859_ _15907_/CLK _15859_/D vssd1 vssd1 vccd1 vccd1 _15859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08400_ _15017_/A _08400_/B _08400_/C vssd1 vssd1 vccd1 vccd1 _08401_/A sky130_fd_sc_hd__and3_1
X_09380_ _15363_/Q _09496_/B _09380_/C vssd1 vssd1 vccd1 vccd1 _09380_/X sky130_fd_sc_hd__and3_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ _08373_/A _08444_/A vssd1 vssd1 vccd1 vccd1 _08331_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_33_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08262_ _08322_/A _08322_/B vssd1 vssd1 vccd1 vccd1 _08263_/B sky130_fd_sc_hd__xor2_4
XFILLER_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08193_ _08193_/A _08291_/A vssd1 vssd1 vccd1 vccd1 _08292_/A sky130_fd_sc_hd__xor2_4
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07977_ _07977_/A _08184_/A vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__xor2_4
XFILLER_68_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09716_ _09748_/C vssd1 vssd1 vccd1 vccd1 _09754_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09647_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _09648_/B sky130_fd_sc_hd__nor2_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _15393_/Q _09585_/C _09404_/X vssd1 vssd1 vccd1 vccd1 _09578_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_70_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08611_/A _08529_/B _08535_/B vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__nor3_1
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11540_ _11826_/A vssd1 vssd1 vccd1 vccd1 _11661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ _15689_/Q _11533_/B _11479_/C vssd1 vssd1 vccd1 vccd1 _11471_/X sky130_fd_sc_hd__and3_1
XFILLER_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10422_ _10444_/A _10422_/B _10422_/C vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__and3_1
X_13210_ _15980_/Q _15979_/Q _15978_/Q _13209_/X vssd1 vssd1 vccd1 vccd1 _15963_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_137_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14190_ _14408_/A vssd1 vssd1 vccd1 vccd1 _14190_/X sky130_fd_sc_hd__clkbuf_2
X_10353_ _10353_/A _10353_/B _10360_/A vssd1 vssd1 vccd1 vccd1 _15513_/D sky130_fd_sc_hd__nor3_1
X_13141_ _13141_/A _13141_/B vssd1 vssd1 vccd1 vccd1 _13142_/B sky130_fd_sc_hd__nor2_1
XFILLER_137_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13072_ _15943_/Q _13078_/C _12855_/X vssd1 vssd1 vccd1 vccd1 _13072_/Y sky130_fd_sc_hd__a21oi_1
X_10284_ _10284_/A _10284_/B _10284_/C vssd1 vssd1 vccd1 vccd1 _10286_/B sky130_fd_sc_hd__or3_1
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12023_ _12055_/C vssd1 vssd1 vccd1 vccd1 _12062_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13974_ _16115_/Q _16114_/Q _16113_/Q _13973_/X vssd1 vssd1 vccd1 vccd1 _16098_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_74_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15713_ _15794_/CLK _15713_/D vssd1 vssd1 vccd1 vccd1 _15713_/Q sky130_fd_sc_hd__dfxtp_1
X_12925_ _12959_/A _12925_/B _12925_/C vssd1 vssd1 vccd1 vccd1 _12926_/A sky130_fd_sc_hd__and3_1
X_15644_ _15655_/CLK _15644_/D vssd1 vssd1 vccd1 vccd1 _15644_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _15906_/Q _12861_/C _12855_/X vssd1 vssd1 vccd1 vccd1 _12856_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11804_/X _11806_/Y _11801_/B _11802_/C vssd1 vssd1 vccd1 vccd1 _11809_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15575_ _15575_/CLK _15575_/D vssd1 vssd1 vccd1 vccd1 _15575_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12784_/X _12785_/Y _12786_/Y _12782_/C vssd1 vssd1 vccd1 vccd1 _12789_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _16214_/Q _14525_/C _07674_/A vssd1 vssd1 vccd1 vccd1 _14527_/B sky130_fd_sc_hd__a21o_1
X_11738_ _11796_/A _11738_/B _11742_/A vssd1 vssd1 vccd1 vccd1 _15729_/D sky130_fd_sc_hd__nor3_1
X_14457_ _14413_/X _14454_/B _14456_/Y vssd1 vssd1 vccd1 vccd1 _16195_/D sky130_fd_sc_hd__o21a_1
X_11669_ _11842_/A vssd1 vssd1 vccd1 vccd1 _11708_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13408_ _13408_/A _13408_/B _13408_/C vssd1 vssd1 vccd1 vccd1 _13410_/B sky130_fd_sc_hd__or3_1
X_14388_ _14388_/A vssd1 vssd1 vccd1 vccd1 _16181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16127_ _16129_/CLK _16127_/D vssd1 vssd1 vccd1 vccd1 _16127_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13339_ _13339_/A _13339_/B _13339_/C vssd1 vssd1 vccd1 vccd1 _13340_/A sky130_fd_sc_hd__and3_1
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16058_ _16060_/CLK _16058_/D vssd1 vssd1 vccd1 vccd1 _16058_/Q sky130_fd_sc_hd__dfxtp_1
X_15009_ _15009_/A _15009_/B vssd1 vssd1 vccd1 vccd1 _16320_/D sky130_fd_sc_hd__nor2_1
X_07900_ _16026_/Q vssd1 vssd1 vccd1 vccd1 _13626_/C sky130_fd_sc_hd__clkinv_4
X_08880_ _15286_/Q _09001_/B _08880_/C vssd1 vssd1 vccd1 vccd1 _08891_/A sky130_fd_sc_hd__and3_1
XFILLER_123_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07831_ _15494_/Q vssd1 vssd1 vccd1 vccd1 _10234_/A sky130_fd_sc_hd__clkinv_2
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07762_ _16278_/Q vssd1 vssd1 vccd1 vccd1 _08099_/A sky130_fd_sc_hd__clkinv_2
X_09501_ _09519_/A _09501_/B _09501_/C vssd1 vssd1 vccd1 vccd1 _09502_/A sky130_fd_sc_hd__and3_1
X_07693_ input7/X vssd1 vssd1 vccd1 vccd1 _10969_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09432_ _15371_/Q _09432_/B _09438_/C vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__nand3_1
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09363_ _09362_/B _09362_/C _09307_/X vssd1 vssd1 vccd1 vccd1 _09364_/C sky130_fd_sc_hd__o21ai_1
XFILLER_80_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08314_ _08315_/A _08315_/B vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__or2_1
X_09294_ _09300_/A _09291_/Y _09293_/Y _09288_/C vssd1 vssd1 vccd1 vccd1 _09296_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_10 _13420_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _15050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 _15972_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ _08246_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _08384_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08176_ _08155_/A _08155_/B _08175_/Y vssd1 vssd1 vccd1 vccd1 _08268_/A sky130_fd_sc_hd__a21o_1
XFILLER_4_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10971_ _15610_/Q _10970_/B _10911_/X vssd1 vssd1 vccd1 vccd1 _10972_/B sky130_fd_sc_hd__a21oi_1
X_12710_ _15883_/Q _12748_/C _12481_/X vssd1 vssd1 vccd1 vccd1 _12712_/B sky130_fd_sc_hd__a21oi_1
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13690_ _13735_/A _13690_/B _13690_/C vssd1 vssd1 vccd1 vccd1 _13691_/A sky130_fd_sc_hd__and3_1
XFILLER_16_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12641_ _12640_/B _12640_/C _12472_/X vssd1 vssd1 vccd1 vccd1 _12642_/C sky130_fd_sc_hd__o21ai_1
X_15360_ _15395_/CLK _15360_/D vssd1 vssd1 vccd1 vccd1 _15360_/Q sky130_fd_sc_hd__dfxtp_2
X_12572_ _12578_/A _12570_/Y _12571_/Y _12565_/C vssd1 vssd1 vccd1 vccd1 _12574_/B
+ sky130_fd_sc_hd__o211a_1
X_14311_ _14308_/A _14308_/B _14307_/Y _14310_/Y vssd1 vssd1 vccd1 vccd1 _16165_/D
+ sky130_fd_sc_hd__o31a_1
X_11523_ _11538_/A _11523_/B _11523_/C vssd1 vssd1 vccd1 vccd1 _11524_/A sky130_fd_sc_hd__and3_1
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15291_ _15301_/CLK _15291_/D vssd1 vssd1 vccd1 vccd1 _15291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14242_ _14242_/A _14242_/B vssd1 vssd1 vccd1 vccd1 _16151_/D sky130_fd_sc_hd__nor2_1
X_11454_ _11454_/A _11454_/B _11454_/C vssd1 vssd1 vccd1 vccd1 _11455_/C sky130_fd_sc_hd__nand3_1
XFILLER_7_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _10577_/A _10405_/B _10405_/C vssd1 vssd1 vccd1 vccd1 _10407_/B sky130_fd_sc_hd__or3_1
X_11385_ _11385_/A vssd1 vssd1 vccd1 vccd1 _15673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14173_ _14179_/A _14172_/Y _14168_/B _14169_/C vssd1 vssd1 vccd1 vccd1 _14175_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13124_ _13122_/Y _13114_/C _13117_/X _13118_/Y vssd1 vssd1 vccd1 vccd1 _13125_/C
+ sky130_fd_sc_hd__a211o_1
X_10336_ _10336_/A _10336_/B vssd1 vssd1 vccd1 vccd1 _10337_/B sky130_fd_sc_hd__nor2_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10267_ _10267_/A vssd1 vssd1 vccd1 vccd1 _15499_/D sky130_fd_sc_hd__clkbuf_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _13069_/A _13055_/B _13055_/C vssd1 vssd1 vccd1 vccd1 _13056_/A sky130_fd_sc_hd__and3_1
XFILLER_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12006_ _12084_/A _12006_/B _12010_/B vssd1 vssd1 vccd1 vccd1 _15770_/D sky130_fd_sc_hd__nor3_1
X_10198_ _15490_/Q _10199_/C _10083_/X vssd1 vssd1 vccd1 vccd1 _10198_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13957_ _16097_/Q _14137_/B _13957_/C vssd1 vssd1 vccd1 vccd1 _13957_/X sky130_fd_sc_hd__and3_1
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12908_ _15915_/Q _13071_/B _12908_/C vssd1 vssd1 vccd1 vccd1 _12917_/A sky130_fd_sc_hd__and3_1
XFILLER_62_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13888_ _13881_/B _13882_/C _13895_/A _13886_/Y vssd1 vssd1 vccd1 vccd1 _13895_/B
+ sky130_fd_sc_hd__a211oi_1
X_15627_ _15194_/Q _15627_/D vssd1 vssd1 vccd1 vccd1 _15627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12839_ _15904_/Q _12840_/C _12668_/X vssd1 vssd1 vccd1 vccd1 _12839_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15558_ _15655_/CLK _15558_/D vssd1 vssd1 vccd1 vccd1 _15558_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14509_ _14510_/B _14510_/C _14510_/A vssd1 vssd1 vccd1 vccd1 _14511_/B sky130_fd_sc_hd__a21o_1
X_15489_ _15224_/Q _15489_/D vssd1 vssd1 vccd1 vccd1 _15489_/Q sky130_fd_sc_hd__dfxtp_1
X_08030_ _15899_/Q _08030_/B vssd1 vssd1 vccd1 vccd1 _08030_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09981_ _11137_/A vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08932_ _08928_/X _08930_/Y _08931_/Y _08924_/C vssd1 vssd1 vccd1 vccd1 _08934_/B
+ sky130_fd_sc_hd__o211ai_1
X_08863_ _08878_/A _08863_/B _08863_/C vssd1 vssd1 vccd1 vccd1 _08864_/A sky130_fd_sc_hd__and3_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07814_ _15755_/Q _15773_/Q vssd1 vssd1 vccd1 vccd1 _07815_/C sky130_fd_sc_hd__or2_1
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08794_ _15272_/Q _08794_/B _08802_/C vssd1 vssd1 vccd1 vccd1 _08799_/A sky130_fd_sc_hd__and3_1
X_07745_ _15413_/Q _08113_/B vssd1 vssd1 vccd1 vccd1 _08107_/B sky130_fd_sc_hd__xnor2_4
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07676_ _14459_/A vssd1 vssd1 vccd1 vccd1 _14648_/A sky130_fd_sc_hd__buf_2
X_09415_ _09415_/A _09415_/B vssd1 vssd1 vccd1 vccd1 _09419_/C sky130_fd_sc_hd__nor2_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09346_ _09346_/A vssd1 vssd1 vccd1 vccd1 _15356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09277_ _15347_/Q _09278_/C _09220_/X vssd1 vssd1 vccd1 vccd1 _09277_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08228_ _08305_/A _08228_/B vssd1 vssd1 vccd1 vccd1 _08228_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08159_ _08159_/A _08174_/A vssd1 vssd1 vccd1 vccd1 _08171_/A sky130_fd_sc_hd__xnor2_4
XFILLER_106_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11170_ _15642_/Q _11178_/C _10940_/X vssd1 vssd1 vccd1 vccd1 _11170_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10121_ _10121_/A vssd1 vssd1 vccd1 vccd1 _10135_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10052_ _10341_/A vssd1 vssd1 vccd1 vccd1 _10284_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14860_ _16292_/Q _14875_/C _14702_/X vssd1 vssd1 vccd1 vccd1 _14862_/B sky130_fd_sc_hd__a21oi_1
XFILLER_87_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13811_ _13809_/A _13809_/B _13810_/X vssd1 vssd1 vccd1 vccd1 _16068_/D sky130_fd_sc_hd__a21oi_1
X_14791_ _14798_/A _14790_/Y _14785_/B _14786_/C vssd1 vssd1 vccd1 vccd1 _14793_/B
+ sky130_fd_sc_hd__o211a_1
X_13742_ _13789_/A _13742_/B _13742_/C vssd1 vssd1 vccd1 vccd1 _13743_/A sky130_fd_sc_hd__and3_1
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10954_ _10954_/A vssd1 vssd1 vccd1 vccd1 _15606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13673_ _13701_/C vssd1 vssd1 vccd1 vccd1 _13707_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_73_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10885_ _10879_/B _10880_/C _10882_/X _10883_/Y vssd1 vssd1 vccd1 vccd1 _10886_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15412_ _15484_/CLK _15412_/D vssd1 vssd1 vccd1 vccd1 _15412_/Q sky130_fd_sc_hd__dfxtp_1
X_12624_ _15870_/Q _12630_/C _12569_/X vssd1 vssd1 vccd1 vccd1 _12624_/Y sky130_fd_sc_hd__a21oi_1
X_15343_ _15348_/CLK _15343_/D vssd1 vssd1 vccd1 vccd1 _15343_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _12552_/X _12553_/Y _12554_/Y _12550_/C vssd1 vssd1 vccd1 vccd1 _12557_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _15694_/Q _11547_/C _11336_/X vssd1 vssd1 vccd1 vccd1 _11509_/B sky130_fd_sc_hd__a21oi_1
X_15274_ _15274_/CLK _15274_/D vssd1 vssd1 vccd1 vccd1 _15274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12486_ _15848_/Q _12492_/C _12370_/X vssd1 vssd1 vccd1 vccd1 _12488_/C sky130_fd_sc_hd__a21o_1
XFILLER_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14225_ _14224_/X _14223_/Y _14042_/X vssd1 vssd1 vccd1 vccd1 _14225_/Y sky130_fd_sc_hd__a21oi_1
X_11437_ _11435_/A _11435_/B _11436_/X vssd1 vssd1 vccd1 vccd1 _15681_/D sky130_fd_sc_hd__a21oi_1
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14156_ _16151_/Q _16150_/Q _16149_/Q _13973_/X vssd1 vssd1 vccd1 vccd1 _16134_/D
+ sky130_fd_sc_hd__o31a_1
X_11368_ _15672_/Q _11374_/C _11137_/X vssd1 vssd1 vccd1 vccd1 _11368_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _13107_/A vssd1 vssd1 vccd1 vccd1 _15947_/D sky130_fd_sc_hd__clkbuf_1
X_10319_ _15509_/Q _10325_/C _10318_/X vssd1 vssd1 vccd1 vccd1 _10319_/Y sky130_fd_sc_hd__a21oi_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14087_ _16122_/Q _14093_/C _13693_/X vssd1 vssd1 vccd1 vccd1 _14087_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11299_ _11296_/X _11297_/Y _11298_/Y _11293_/C vssd1 vssd1 vccd1 vccd1 _11301_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13051_/C vssd1 vssd1 vccd1 vccd1 _13059_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14989_ hold5/X _14994_/C _14988_/X vssd1 vssd1 vccd1 vccd1 _14989_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09200_ _15335_/Q _09242_/C _09029_/X vssd1 vssd1 vccd1 vccd1 _09202_/B sky130_fd_sc_hd__a21oi_1
XFILLER_22_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09131_ _09129_/A _09129_/B _09130_/X vssd1 vssd1 vccd1 vccd1 _15322_/D sky130_fd_sc_hd__a21oi_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09062_ _15313_/Q _09067_/C _08824_/X vssd1 vssd1 vccd1 vccd1 _09062_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08013_ _14022_/C _07868_/B _08012_/X vssd1 vssd1 vccd1 vccd1 _08014_/B sky130_fd_sc_hd__o21a_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09964_ _15454_/Q _10022_/B _09967_/C vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__and3_1
XFILLER_103_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08915_ _08916_/B _08916_/C _08916_/A vssd1 vssd1 vccd1 vccd1 _08917_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09895_ _15442_/Q _09950_/B _09903_/C vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__and3_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _08867_/C vssd1 vssd1 vccd1 vccd1 _08880_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08777_ _08783_/B _08777_/B vssd1 vssd1 vccd1 vccd1 _08779_/A sky130_fd_sc_hd__or2_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07728_ _09367_/A _07728_/B vssd1 vssd1 vccd1 vccd1 _07729_/B sky130_fd_sc_hd__xnor2_2
XFILLER_25_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07659_ input4/X vssd1 vssd1 vccd1 vccd1 _10947_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10670_ _11303_/A vssd1 vssd1 vccd1 vccd1 _10895_/B sky130_fd_sc_hd__buf_2
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _09323_/B _09324_/C _09326_/X _09327_/Y vssd1 vssd1 vccd1 vccd1 _09330_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _15825_/Q _12346_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12340_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12271_ _12268_/X _12269_/Y _12270_/Y _12266_/C vssd1 vssd1 vccd1 vccd1 _12273_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_5_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _15186_/A _14010_/B vssd1 vssd1 vccd1 vccd1 _14011_/B sky130_fd_sc_hd__and2_1
X_11222_ _11222_/A vssd1 vssd1 vccd1 vccd1 _11222_/X sky130_fd_sc_hd__buf_2
XFILLER_141_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _11189_/A _11153_/B _11153_/C vssd1 vssd1 vccd1 vccd1 _11154_/A sky130_fd_sc_hd__and3_1
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10104_ _10102_/Y _10097_/C _10109_/A _10101_/Y vssd1 vssd1 vccd1 vccd1 _10109_/B
+ sky130_fd_sc_hd__a211oi_1
X_11084_ _11082_/Y _11076_/C _11089_/A _11079_/Y vssd1 vssd1 vccd1 vccd1 _11089_/B
+ sky130_fd_sc_hd__a211oi_1
X_15961_ _15961_/CLK _15961_/D vssd1 vssd1 vccd1 vccd1 _15961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10035_ _10035_/A _10035_/B _10035_/C vssd1 vssd1 vccd1 vccd1 _10036_/A sky130_fd_sc_hd__and3_1
XFILLER_88_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14912_ _16303_/Q _14916_/C _14789_/X vssd1 vssd1 vccd1 vccd1 _14912_/Y sky130_fd_sc_hd__a21oi_1
X_15892_ _15907_/CLK _15892_/D vssd1 vssd1 vccd1 vccd1 _15892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14843_ _14843_/A _14843_/B vssd1 vssd1 vccd1 vccd1 _14843_/X sky130_fd_sc_hd__or2_1
XFILLER_64_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14774_ _07707_/X _14771_/A _14773_/Y vssd1 vssd1 vccd1 vccd1 _16268_/D sky130_fd_sc_hd__o21a_1
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11986_ _15768_/Q _11986_/B _11986_/C vssd1 vssd1 vccd1 vccd1 _11986_/Y sky130_fd_sc_hd__nand3_1
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13725_ _13729_/C vssd1 vssd1 vccd1 vccd1 _13738_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10937_ _10960_/A _10937_/B _10937_/C vssd1 vssd1 vccd1 vccd1 _10938_/A sky130_fd_sc_hd__and3_1
XFILLER_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13656_ _16043_/Q _13655_/C _13452_/X vssd1 vssd1 vccd1 vccd1 _13657_/B sky130_fd_sc_hd__a21oi_1
X_10868_ _15593_/Q vssd1 vssd1 vccd1 vccd1 _10882_/C sky130_fd_sc_hd__clkinv_2
XFILLER_32_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12607_ _15868_/Q _12667_/B _12610_/C vssd1 vssd1 vccd1 vccd1 _12607_/X sky130_fd_sc_hd__and3_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13587_ _13595_/A _13587_/B _13587_/C vssd1 vssd1 vccd1 vccd1 _13588_/A sky130_fd_sc_hd__and3_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _15583_/Q _10798_/C _10624_/X vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__a21oi_1
XFILLER_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15326_ _15333_/CLK _15326_/D vssd1 vssd1 vccd1 vccd1 _15326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12538_ _15856_/Q _12593_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12543_/A sky130_fd_sc_hd__and3_1
XFILLER_118_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15257_ _15274_/CLK _15257_/D vssd1 vssd1 vccd1 vccd1 _15257_/Q sky130_fd_sc_hd__dfxtp_1
X_12469_ _13029_/A vssd1 vssd1 vccd1 vccd1 _12698_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14208_ _14208_/A _14208_/B _14212_/A vssd1 vssd1 vccd1 vccd1 _16144_/D sky130_fd_sc_hd__nor3_1
XFILLER_125_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15188_ _15188_/A _15188_/B vssd1 vssd1 vccd1 vccd1 _16365_/D sky130_fd_sc_hd__nor2_1
XFILLER_141_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14139_ _14137_/X _14139_/B vssd1 vssd1 vccd1 vccd1 _14139_/X sky130_fd_sc_hd__and2b_1
XFILLER_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08700_ _15258_/Q _08706_/C _08575_/X vssd1 vssd1 vccd1 vccd1 _08700_/Y sky130_fd_sc_hd__a21oi_1
X_09680_ _15408_/Q _09911_/B _09680_/C vssd1 vssd1 vccd1 vccd1 _09680_/Y sky130_fd_sc_hd__nand3_1
X_08631_ _12668_/A vssd1 vssd1 vccd1 vccd1 _08865_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08562_ _08560_/X _08561_/Y _08557_/B _08558_/C vssd1 vssd1 vccd1 vccd1 _08564_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08493_ _15229_/Q _10939_/C _08493_/C vssd1 vssd1 vccd1 vccd1 _08493_/X sky130_fd_sc_hd__and3_1
XFILLER_23_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09114_ _09112_/Y _09108_/C _09110_/X _09111_/Y vssd1 vssd1 vccd1 vccd1 _09115_/C
+ sky130_fd_sc_hd__a211o_1
X_09045_ _15311_/Q _09158_/B _09047_/C vssd1 vssd1 vccd1 vccd1 _09045_/X sky130_fd_sc_hd__and3_1
XFILLER_117_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09947_ _09967_/C vssd1 vssd1 vccd1 vccd1 _09979_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09878_ _09878_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _09883_/C sky130_fd_sc_hd__nor2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08829_ _08909_/A _08829_/B _08834_/B vssd1 vssd1 vccd1 vccd1 _15276_/D sky130_fd_sc_hd__nor3_1
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11840_ _12068_/A _11843_/C vssd1 vssd1 vccd1 vccd1 _11840_/X sky130_fd_sc_hd__or2_1
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11769_/Y _11765_/C _11778_/A _11768_/Y vssd1 vssd1 vccd1 vccd1 _11778_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _13713_/A _13512_/C vssd1 vssd1 vccd1 vccd1 _13510_/X sky130_fd_sc_hd__or2_1
X_10722_ _15570_/Q _10778_/B _10722_/C vssd1 vssd1 vccd1 vccd1 _10722_/Y sky130_fd_sc_hd__nand3_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _14485_/Y _14488_/X _14489_/Y vssd1 vssd1 vccd1 vccd1 _16202_/D sky130_fd_sc_hd__o21a_1
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ _13439_/Y _13434_/C _13436_/X _13438_/Y vssd1 vssd1 vccd1 vccd1 _13442_/C
+ sky130_fd_sc_hd__a211o_1
X_10653_ _10653_/A vssd1 vssd1 vccd1 vccd1 _15559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16160_ _16187_/CLK _16160_/D vssd1 vssd1 vccd1 vccd1 _16160_/Q sky130_fd_sc_hd__dfxtp_1
X_13372_ _15993_/Q _13420_/B _13372_/C vssd1 vssd1 vccd1 vccd1 _13377_/A sky130_fd_sc_hd__and3_1
XFILLER_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ _10604_/C vssd1 vssd1 vccd1 vccd1 _10617_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15111_ _15111_/A _15111_/B vssd1 vssd1 vccd1 vccd1 _15112_/B sky130_fd_sc_hd__nor2_1
X_12323_ _15823_/Q _12383_/B _12326_/C vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__and3_1
X_16091_ _16224_/CLK _16091_/D vssd1 vssd1 vccd1 vccd1 _16091_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15042_ _15040_/A _15040_/B _15041_/X vssd1 vssd1 vccd1 vccd1 _16327_/D sky130_fd_sc_hd__a21oi_1
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12254_ _15811_/Q _12309_/B _12262_/C vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__and3_1
XFILLER_141_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11205_ _11203_/A _11203_/B _11204_/X vssd1 vssd1 vccd1 vccd1 _15645_/D sky130_fd_sc_hd__a21oi_1
XFILLER_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ _13029_/A vssd1 vssd1 vccd1 vccd1 _12413_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11136_ _15636_/Q _11367_/B _11136_/C vssd1 vssd1 vccd1 vccd1 _11146_/A sky130_fd_sc_hd__and3_1
XFILLER_110_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11067_ _11064_/X _11065_/Y _11066_/Y _11062_/C vssd1 vssd1 vccd1 vccd1 _11069_/B
+ sky130_fd_sc_hd__o211ai_1
X_15944_ _15196_/Q _15944_/D vssd1 vssd1 vccd1 vccd1 _15944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10018_ _10016_/X _10017_/Y _10013_/B _10014_/C vssd1 vssd1 vccd1 vccd1 _10020_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15875_ _07603_/A _15875_/D vssd1 vssd1 vccd1 vccd1 _15875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14826_ _16284_/Q _14941_/B _14826_/C vssd1 vssd1 vccd1 vccd1 _14829_/B sky130_fd_sc_hd__nand3_1
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14757_ _14757_/A _14757_/B vssd1 vssd1 vccd1 vccd1 _14759_/A sky130_fd_sc_hd__or2_1
XFILLER_44_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11969_ _15766_/Q _12007_/C _11912_/X vssd1 vssd1 vccd1 vccd1 _11971_/B sky130_fd_sc_hd__a21oi_1
XFILLER_44_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13708_ _14099_/B vssd1 vssd1 vccd1 vccd1 _13708_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14688_ _07675_/X _14679_/A _14683_/B _14687_/Y vssd1 vssd1 vccd1 vccd1 _16247_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_32_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13639_ _13639_/A vssd1 vssd1 vccd1 vccd1 _16038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16358_ _16358_/CLK _16358_/D vssd1 vssd1 vccd1 vccd1 _16358_/Q sky130_fd_sc_hd__dfxtp_1
X_15309_ _15333_/CLK _15309_/D vssd1 vssd1 vccd1 vccd1 _15309_/Q sky130_fd_sc_hd__dfxtp_1
X_16289_ _16304_/CLK _16289_/D vssd1 vssd1 vccd1 vccd1 _16289_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09801_ _09801_/A vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07993_ _14584_/C _07874_/B _07873_/B vssd1 vssd1 vccd1 vccd1 _07999_/A sky130_fd_sc_hd__o21ai_1
XFILLER_87_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09732_ _09732_/A vssd1 vssd1 vccd1 vccd1 _15416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09663_ _15406_/Q _09663_/B _09671_/C vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__and3_1
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08614_ _15246_/Q _08853_/B _08622_/C vssd1 vssd1 vccd1 vccd1 _08619_/B sky130_fd_sc_hd__nand3_1
XFILLER_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09594_ _09708_/A _09594_/B _09594_/C vssd1 vssd1 vccd1 vccd1 _09598_/B sky130_fd_sc_hd__or3_1
XFILLER_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08545_ _15251_/Q _15250_/Q _15249_/Q _07608_/X vssd1 vssd1 vccd1 vccd1 _15234_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _08505_/C vssd1 vssd1 vccd1 vccd1 _08522_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09028_ _14901_/A vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__buf_4
XFILLER_2_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13990_ _16104_/Q _14988_/A _13990_/C vssd1 vssd1 vccd1 vccd1 _13998_/A sky130_fd_sc_hd__and3_1
XFILLER_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _15921_/Q _12996_/B _12941_/C vssd1 vssd1 vccd1 vccd1 _12941_/X sky130_fd_sc_hd__and3_1
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15660_ _15763_/CLK _15660_/D vssd1 vssd1 vccd1 vccd1 _15660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12872_ _12872_/A vssd1 vssd1 vccd1 vccd1 _15907_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14806_/A _14611_/B vssd1 vssd1 vccd1 vccd1 _14612_/B sky130_fd_sc_hd__and2_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _11821_/Y _11817_/C _11819_/X _11820_/Y vssd1 vssd1 vccd1 vccd1 _11824_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15591_ _15194_/Q _15591_/D vssd1 vssd1 vccd1 vccd1 _15591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14936_/A vssd1 vssd1 vccd1 vccd1 _14626_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _15732_/Q _11986_/B _11754_/C vssd1 vssd1 vccd1 vccd1 _11754_/Y sky130_fd_sc_hd__nand3_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _15568_/Q _10817_/B _10714_/C vssd1 vssd1 vccd1 vccd1 _10710_/A sky130_fd_sc_hd__and3_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14473_/A vssd1 vssd1 vccd1 vccd1 _16199_/D sky130_fd_sc_hd__clkbuf_1
X_11685_ _11686_/B _11686_/C _11686_/A vssd1 vssd1 vccd1 vccd1 _11687_/B sky130_fd_sc_hd__a21o_1
XFILLER_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16212_ _16222_/CLK _16212_/D vssd1 vssd1 vccd1 vccd1 _16212_/Q sky130_fd_sc_hd__dfxtp_1
X_13424_ _16003_/Q _13628_/B _13430_/C vssd1 vssd1 vccd1 vccd1 _13427_/B sky130_fd_sc_hd__nand3_1
X_10636_ _10676_/A _10636_/B _10636_/C vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__and3_1
XFILLER_127_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16143_ _16143_/CLK _16143_/D vssd1 vssd1 vccd1 vccd1 _16143_/Q sky130_fd_sc_hd__dfxtp_1
X_13355_ _13353_/A _13353_/B _13354_/X vssd1 vssd1 vccd1 vccd1 _15987_/D sky130_fd_sc_hd__a21oi_1
X_10567_ _10645_/A _10567_/B _10572_/B vssd1 vssd1 vccd1 vccd1 _15545_/D sky130_fd_sc_hd__nor3_1
XFILLER_6_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12306_ _12326_/C vssd1 vssd1 vccd1 vccd1 _12339_/C sky130_fd_sc_hd__clkbuf_1
X_16074_ _16143_/CLK _16074_/D vssd1 vssd1 vccd1 vccd1 _16074_/Q sky130_fd_sc_hd__dfxtp_1
X_13286_ _15977_/Q _13286_/B _13291_/C vssd1 vssd1 vccd1 vccd1 _13286_/Y sky130_fd_sc_hd__nand3_1
X_10498_ _15536_/Q _10506_/C _10318_/X vssd1 vssd1 vccd1 vccd1 _10498_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15025_ _16329_/Q _15024_/C _14942_/X vssd1 vssd1 vccd1 vccd1 _15027_/C sky130_fd_sc_hd__a21o_1
X_12237_ _12243_/B _12237_/B vssd1 vssd1 vccd1 vccd1 _12239_/A sky130_fd_sc_hd__or2_1
XFILLER_142_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12168_ _12165_/X _12166_/Y _12167_/Y _12162_/C vssd1 vssd1 vccd1 vccd1 _12170_/B
+ sky130_fd_sc_hd__o211ai_1
X_11119_ _15634_/Q _11236_/B _11121_/C vssd1 vssd1 vccd1 vccd1 _11119_/X sky130_fd_sc_hd__and3_1
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12099_ _15787_/Q _12099_/B _12102_/C vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__and3_1
XFILLER_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 in1[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_6
X_15927_ _15196_/Q _15927_/D vssd1 vssd1 vccd1 vccd1 _15927_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15858_ _15907_/CLK _15858_/D vssd1 vssd1 vccd1 vccd1 _15858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14809_ _14766_/X _14811_/C _14808_/X vssd1 vssd1 vccd1 vccd1 _14810_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15789_ _15195_/Q _15789_/D vssd1 vssd1 vccd1 vccd1 _15789_/Q sky130_fd_sc_hd__dfxtp_1
X_08330_ _08330_/A _08330_/B vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__xnor2_4
XFILLER_33_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08261_ _08147_/A _08147_/B _08260_/Y vssd1 vssd1 vccd1 vccd1 _08322_/B sky130_fd_sc_hd__a21oi_2
X_08192_ _08295_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08291_/A sky130_fd_sc_hd__nand2_2
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07976_ _07976_/A _07976_/B vssd1 vssd1 vccd1 vccd1 _08184_/A sky130_fd_sc_hd__xnor2_2
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09715_ _09735_/C vssd1 vssd1 vccd1 vccd1 _09748_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09646_ _09652_/B _09646_/B vssd1 vssd1 vccd1 vccd1 _09648_/A sky130_fd_sc_hd__or2_1
XFILLER_16_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09577_ _15393_/Q _09577_/B _09577_/C vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__and3_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _08526_/Y _08519_/C _08535_/A _08525_/Y vssd1 vssd1 vccd1 vccd1 _08535_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08459_ _14163_/A vssd1 vssd1 vccd1 vccd1 _13972_/A sky130_fd_sc_hd__clkbuf_2
X_11470_ _11470_/A vssd1 vssd1 vccd1 vccd1 _15687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10421_ _10421_/A _10421_/B _10421_/C vssd1 vssd1 vccd1 vccd1 _10422_/C sky130_fd_sc_hd__nand3_1
XFILLER_136_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13140_ _13146_/B _13140_/B vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__or2_1
X_10352_ _15514_/Q _10532_/B _10363_/C vssd1 vssd1 vccd1 vccd1 _10360_/A sky130_fd_sc_hd__and3_1
X_13071_ _15943_/Q _13071_/B _13071_/C vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__and3_1
X_10283_ _10404_/A vssd1 vssd1 vccd1 vccd1 _10323_/A sky130_fd_sc_hd__clkbuf_2
X_12022_ _12042_/C vssd1 vssd1 vccd1 vccd1 _12055_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_78_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13973_ _14818_/A vssd1 vssd1 vccd1 vccd1 _13973_/X sky130_fd_sc_hd__buf_2
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15712_ _15794_/CLK _15712_/D vssd1 vssd1 vccd1 vccd1 _15712_/Q sky130_fd_sc_hd__dfxtp_1
X_12924_ _12923_/B _12923_/C _12758_/X vssd1 vssd1 vccd1 vccd1 _12925_/C sky130_fd_sc_hd__o21ai_1
XFILLER_74_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15643_ _15194_/Q _15643_/D vssd1 vssd1 vccd1 vccd1 _15643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12855_ _13654_/A vssd1 vssd1 vccd1 vccd1 _12855_/X sky130_fd_sc_hd__buf_2
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _15741_/Q _11814_/C _11805_/X vssd1 vssd1 vccd1 vccd1 _11806_/Y sky130_fd_sc_hd__a21oi_1
X_15574_ _15655_/CLK _15574_/D vssd1 vssd1 vccd1 vccd1 _15574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _15894_/Q _12840_/B _12786_/C vssd1 vssd1 vccd1 vccd1 _12786_/Y sky130_fd_sc_hd__nand3_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _16214_/Q _14566_/B _14525_/C vssd1 vssd1 vccd1 vccd1 _14525_/X sky130_fd_sc_hd__and3_1
X_11737_ _15730_/Q _11737_/B _11745_/C vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__and3_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14456_ _14368_/X _14454_/B _14415_/X vssd1 vssd1 vccd1 vccd1 _14456_/Y sky130_fd_sc_hd__a21oi_1
X_11668_ _11666_/A _11666_/B _11667_/X vssd1 vssd1 vccd1 vccd1 _15717_/D sky130_fd_sc_hd__a21oi_1
X_13407_ _13405_/A _13405_/B _13406_/X vssd1 vssd1 vccd1 vccd1 _15996_/D sky130_fd_sc_hd__a21oi_1
X_10619_ _15554_/Q _10681_/B _10623_/C vssd1 vssd1 vccd1 vccd1 _10619_/Y sky130_fd_sc_hd__nand3_1
X_14387_ _14552_/A _14387_/B _14387_/C vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__and3_1
X_11599_ _15708_/Q _11655_/B _11599_/C vssd1 vssd1 vccd1 vccd1 _11608_/A sky130_fd_sc_hd__and3_1
X_16126_ _16129_/CLK _16126_/D vssd1 vssd1 vccd1 vccd1 _16126_/Q sky130_fd_sc_hd__dfxtp_2
X_13338_ _13336_/Y _13331_/C _13333_/X _13334_/Y vssd1 vssd1 vccd1 vccd1 _13339_/C
+ sky130_fd_sc_hd__a211o_1
X_16057_ _16060_/CLK _16057_/D vssd1 vssd1 vccd1 vccd1 _16057_/Q sky130_fd_sc_hd__dfxtp_1
X_13269_ _13526_/A vssd1 vssd1 vccd1 vccd1 _13269_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15008_ _14964_/X _15010_/C _15007_/X vssd1 vssd1 vccd1 vccd1 _15009_/B sky130_fd_sc_hd__o21ai_1
X_07830_ _15404_/Q vssd1 vssd1 vccd1 vccd1 _09658_/A sky130_fd_sc_hd__inv_2
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ _16260_/Q vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__clkinv_2
XFILLER_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09500_ _09493_/B _09494_/C _09496_/X _09498_/Y vssd1 vssd1 vccd1 vccd1 _09501_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07692_ _07692_/A _07692_/B vssd1 vssd1 vccd1 vccd1 _15203_/D sky130_fd_sc_hd__nor2_1
XFILLER_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09431_ _09487_/A _09431_/B _09435_/A vssd1 vssd1 vccd1 vccd1 _15369_/D sky130_fd_sc_hd__nor3_1
XFILLER_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ _09419_/A _09362_/B _09362_/C vssd1 vssd1 vccd1 vccd1 _09364_/B sky130_fd_sc_hd__or3_1
XFILLER_33_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08313_ _08255_/A _08255_/B _08312_/Y vssd1 vssd1 vccd1 vccd1 _08315_/B sky130_fd_sc_hd__a21oi_1
X_09293_ _15348_/Q _09524_/B _09297_/C vssd1 vssd1 vccd1 vccd1 _09293_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_11 _11080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _13919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_33 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ _08244_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _08246_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08175_ _08175_/A _08175_/B vssd1 vssd1 vccd1 vccd1 _08175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07959_ _12077_/A _07861_/B _07860_/A vssd1 vssd1 vccd1 vccd1 _07976_/A sky130_fd_sc_hd__o21a_2
XFILLER_87_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10970_ _15610_/Q _10970_/B _10970_/C vssd1 vssd1 vccd1 vccd1 _10979_/B sky130_fd_sc_hd__and3_1
XFILLER_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09629_ _15401_/Q _09638_/C _09453_/X vssd1 vssd1 vccd1 vccd1 _09629_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ _12869_/A _12640_/B _12640_/C vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__or3_1
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12571_ _15860_/Q _12744_/B _12575_/C vssd1 vssd1 vccd1 vccd1 _12571_/Y sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_50_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16268_/CLK sky130_fd_sc_hd__clkbuf_16
X_14310_ _14308_/X _14307_/Y _14309_/X vssd1 vssd1 vccd1 vccd1 _14310_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _11515_/B _11516_/C _11518_/X _11520_/Y vssd1 vssd1 vccd1 vccd1 _11523_/C
+ sky130_fd_sc_hd__a211o_1
X_15290_ _15301_/CLK _15290_/D vssd1 vssd1 vccd1 vccd1 _15290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _14061_/X _14153_/X _14235_/B _14240_/X vssd1 vssd1 vccd1 vccd1 _14242_/B
+ sky130_fd_sc_hd__a31o_1
X_11453_ _11454_/B _11454_/C _11454_/A vssd1 vssd1 vccd1 vccd1 _11455_/B sky130_fd_sc_hd__a21o_1
X_10404_ _10404_/A vssd1 vssd1 vccd1 vccd1 _10444_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14172_ _16140_/Q _14171_/C _14033_/X vssd1 vssd1 vccd1 vccd1 _14172_/Y sky130_fd_sc_hd__a21oi_1
X_11384_ _11420_/A _11384_/B _11384_/C vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__and3_1
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13123_ _13117_/X _13118_/Y _13122_/Y _13114_/C vssd1 vssd1 vccd1 vccd1 _13125_/B
+ sky130_fd_sc_hd__o211ai_1
X_10335_ _10342_/B _10335_/B vssd1 vssd1 vccd1 vccd1 _10337_/A sky130_fd_sc_hd__or2_1
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _13048_/B _13049_/C _13051_/X _13052_/Y vssd1 vssd1 vccd1 vccd1 _13055_/C
+ sky130_fd_sc_hd__a211o_1
X_10266_ _10266_/A _10266_/B _10266_/C vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__and3_1
XFILLER_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ _12003_/Y _11997_/C _12010_/A _12002_/Y vssd1 vssd1 vccd1 vccd1 _12010_/B
+ sky130_fd_sc_hd__a211oi_1
X_10197_ _15490_/Q _10310_/B _10199_/C vssd1 vssd1 vccd1 vccd1 _10197_/X sky130_fd_sc_hd__and3_1
XFILLER_87_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13956_ _13953_/B _13952_/Y _13953_/A vssd1 vssd1 vccd1 vccd1 _13956_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_62_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12907_ _12907_/A vssd1 vssd1 vccd1 vccd1 _15913_/D sky130_fd_sc_hd__clkbuf_1
X_13887_ _13895_/A _13886_/Y _13881_/B _13882_/C vssd1 vssd1 vccd1 vccd1 _13889_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15626_ _15194_/Q _15626_/D vssd1 vssd1 vccd1 vccd1 _15626_/Q sky130_fd_sc_hd__dfxtp_1
X_12838_ _15904_/Q _12947_/B _12840_/C vssd1 vssd1 vccd1 vccd1 _12838_/X sky130_fd_sc_hd__and3_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15557_ _15584_/CLK _15557_/D vssd1 vssd1 vccd1 vccd1 _15557_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _15892_/Q _12879_/B _12778_/C vssd1 vssd1 vccd1 vccd1 _12774_/A sky130_fd_sc_hd__and3_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16166_/CLK sky130_fd_sc_hd__clkbuf_16
X_14508_ _16211_/Q _14513_/C _07632_/A vssd1 vssd1 vccd1 vccd1 _14510_/C sky130_fd_sc_hd__a21o_1
XFILLER_148_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15488_ _15224_/Q _15488_/D vssd1 vssd1 vccd1 vccd1 _15488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14439_ _14517_/A _14439_/B _14442_/B vssd1 vssd1 vccd1 vccd1 _16191_/D sky130_fd_sc_hd__nor3_1
XFILLER_116_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16109_ _16119_/CLK _16109_/D vssd1 vssd1 vccd1 vccd1 _16109_/Q sky130_fd_sc_hd__dfxtp_2
X_09980_ _11424_/A vssd1 vssd1 vccd1 vccd1 _11137_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_143_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08931_ _15292_/Q _09047_/B _08931_/C vssd1 vssd1 vccd1 vccd1 _08931_/Y sky130_fd_sc_hd__nand3_1
XFILLER_143_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08862_ _08856_/B _08857_/C _08859_/X _08860_/Y vssd1 vssd1 vccd1 vccd1 _08863_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07813_ _15755_/Q _15773_/Q vssd1 vssd1 vccd1 vccd1 _08052_/A sky130_fd_sc_hd__nand2_1
X_08793_ _15272_/Q _08831_/C _08735_/X vssd1 vssd1 vccd1 vccd1 _08795_/B sky130_fd_sc_hd__a21oi_1
XFILLER_85_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07744_ _15395_/Q _15377_/Q vssd1 vssd1 vccd1 vccd1 _08113_/B sky130_fd_sc_hd__xor2_4
XFILLER_84_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07675_ _15001_/A vssd1 vssd1 vccd1 vccd1 _07675_/X sky130_fd_sc_hd__buf_2
XFILLER_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09414_ _09414_/A _09414_/B vssd1 vssd1 vccd1 vccd1 _09415_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09345_ _09345_/A _09345_/B _09345_/C vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_32_clk clkbuf_opt_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _16242_/CLK sky130_fd_sc_hd__clkbuf_16
X_09276_ _15347_/Q _09444_/B _09278_/C vssd1 vssd1 vccd1 vccd1 _09276_/X sky130_fd_sc_hd__and3_1
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08227_ _08305_/B _08227_/B vssd1 vssd1 vccd1 vccd1 _08228_/B sky130_fd_sc_hd__and2b_1
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08158_ _08173_/A _08173_/B vssd1 vssd1 vccd1 vccd1 _08174_/A sky130_fd_sc_hd__xnor2_2
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08089_ _10639_/A _10527_/A _08088_/Y vssd1 vssd1 vccd1 vccd1 _08103_/A sky130_fd_sc_hd__o21ai_4
X_10120_ _15484_/Q _15483_/Q _15482_/Q _10119_/X vssd1 vssd1 vccd1 vccd1 _15476_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_clk _15665_/CLK vssd1 vssd1 vccd1 vccd1 _15683_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10051_ _10114_/A vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13810_ _14644_/A _13812_/C vssd1 vssd1 vccd1 vccd1 _13810_/X sky130_fd_sc_hd__or2_1
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14790_ hold14/A _14795_/C _14789_/X vssd1 vssd1 vccd1 vccd1 _14790_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13741_ _13734_/B _13735_/C _13738_/X _13739_/Y vssd1 vssd1 vccd1 vccd1 _13742_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10953_ _10960_/A _10953_/B _10953_/C vssd1 vssd1 vccd1 vccd1 _10954_/A sky130_fd_sc_hd__and3_1
XFILLER_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13672_ _13686_/C vssd1 vssd1 vccd1 vccd1 _13701_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10884_ _10882_/X _10883_/Y _10879_/B _10880_/C vssd1 vssd1 vccd1 vccd1 _10886_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15411_ _15484_/CLK _15411_/D vssd1 vssd1 vccd1 vccd1 _15411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12623_ _15870_/Q _12798_/B _12623_/C vssd1 vssd1 vccd1 vccd1 _12634_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_23_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _16148_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15342_ _15359_/CLK _15342_/D vssd1 vssd1 vccd1 vccd1 _15342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12554_ _15858_/Q _12554_/B _12554_/C vssd1 vssd1 vccd1 vccd1 _12554_/Y sky130_fd_sc_hd__nand3_1
X_11505_ _11541_/C vssd1 vssd1 vccd1 vccd1 _11547_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15273_ _15282_/CLK _15273_/D vssd1 vssd1 vccd1 vccd1 _15273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12485_ _15848_/Q _12653_/B _12492_/C vssd1 vssd1 vccd1 vccd1 _12488_/B sky130_fd_sc_hd__nand3_1
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14224_ _14224_/A _14224_/B vssd1 vssd1 vccd1 vccd1 _14224_/X sky130_fd_sc_hd__or2_1
XFILLER_8_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11436_ _11493_/A _11439_/C vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__or2_1
XFILLER_125_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14155_ _14155_/A _14155_/B vssd1 vssd1 vccd1 vccd1 _16133_/D sky130_fd_sc_hd__nor2_1
X_11367_ _15672_/Q _11367_/B _11367_/C vssd1 vssd1 vccd1 vccd1 _11377_/A sky130_fd_sc_hd__and3_1
X_13106_ _13149_/A _13106_/B _13106_/C vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__and3_1
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ _10610_/A vssd1 vssd1 vccd1 vccd1 _10318_/X sky130_fd_sc_hd__clkbuf_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14086_ _16122_/Q _14993_/A _14093_/C vssd1 vssd1 vccd1 vccd1 _14086_/X sky130_fd_sc_hd__and3_1
X_11298_ _15660_/Q _11409_/B _11298_/C vssd1 vssd1 vccd1 vccd1 _11298_/Y sky130_fd_sc_hd__nand3_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _15935_/Q vssd1 vssd1 vccd1 vccd1 _13051_/C sky130_fd_sc_hd__inv_2
X_10249_ _10247_/X _10248_/Y _10244_/B _10245_/C vssd1 vssd1 vccd1 vccd1 _10251_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_79_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14988_ _14988_/A vssd1 vssd1 vccd1 vccd1 _14988_/X sky130_fd_sc_hd__buf_2
XFILLER_75_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ _16094_/Q _13981_/B _13945_/C vssd1 vssd1 vccd1 vccd1 _13942_/B sky130_fd_sc_hd__nand3_1
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _15194_/Q _15609_/D vssd1 vssd1 vccd1 vccd1 _15609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _16022_/CLK sky130_fd_sc_hd__clkbuf_16
X_09130_ _09185_/A _09133_/C vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__or2_1
XFILLER_147_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09061_ _15313_/Q _09290_/B _09061_/C vssd1 vssd1 vccd1 vccd1 _09070_/A sky130_fd_sc_hd__and3_1
X_08012_ _14117_/C _08012_/B vssd1 vssd1 vccd1 vccd1 _08012_/X sky130_fd_sc_hd__or2_1
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09963_ _09963_/A vssd1 vssd1 vccd1 vccd1 _15452_/D sky130_fd_sc_hd__clkbuf_1
X_08914_ _15291_/Q _08919_/C _08913_/X vssd1 vssd1 vccd1 vccd1 _08916_/C sky130_fd_sc_hd__a21o_1
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09894_ _15442_/Q _09931_/C _09893_/X vssd1 vssd1 vccd1 vccd1 _09896_/B sky130_fd_sc_hd__a21oi_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08859_/C vssd1 vssd1 vccd1 vccd1 _08867_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08776_ _15269_/Q _08775_/C _08590_/X vssd1 vssd1 vccd1 vccd1 _08777_/B sky130_fd_sc_hd__a21oi_1
XFILLER_38_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07727_ _07727_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07728_/B sky130_fd_sc_hd__nand2_2
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07658_ _15205_/Q _14755_/B _07658_/C vssd1 vssd1 vccd1 vccd1 _07665_/A sky130_fd_sc_hd__and3_1
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09328_ _09326_/X _09327_/Y _09323_/B _09324_/C vssd1 vssd1 vccd1 vccd1 _09330_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ _09290_/C vssd1 vssd1 vccd1 vccd1 _09297_/C sky130_fd_sc_hd__clkbuf_2
X_12270_ _15813_/Q _12270_/B _12270_/C vssd1 vssd1 vccd1 vccd1 _12270_/Y sky130_fd_sc_hd__nand3_1
XFILLER_107_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11221_ _15650_/Q _11221_/B _11228_/C vssd1 vssd1 vccd1 vccd1 _11225_/B sky130_fd_sc_hd__nand3_1
XFILLER_134_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11152_ _11151_/B _11151_/C _11038_/X vssd1 vssd1 vccd1 vccd1 _11153_/C sky130_fd_sc_hd__o21ai_1
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10103_ _10109_/A _10101_/Y _10102_/Y _10097_/C vssd1 vssd1 vccd1 vccd1 _10105_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11083_ _11089_/A _11079_/Y _11082_/Y _11076_/C vssd1 vssd1 vccd1 vccd1 _11085_/B
+ sky130_fd_sc_hd__o211a_1
X_15960_ _15961_/CLK _15960_/D vssd1 vssd1 vccd1 vccd1 _15960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10034_ _10032_/Y _10027_/C _10029_/X _10031_/Y vssd1 vssd1 vccd1 vccd1 _10035_/C
+ sky130_fd_sc_hd__a211o_1
X_14911_ _16303_/Q _15031_/B _14916_/C vssd1 vssd1 vccd1 vccd1 _14920_/A sky130_fd_sc_hd__and3_1
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15891_ _15907_/CLK _15891_/D vssd1 vssd1 vccd1 vccd1 _15891_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14842_ _14842_/A _14842_/B vssd1 vssd1 vccd1 vccd1 _14843_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11985_ _15769_/Q _11986_/C _11812_/X vssd1 vssd1 vccd1 vccd1 _11985_/Y sky130_fd_sc_hd__a21oi_1
X_14773_ _14772_/X _14771_/A _14614_/X vssd1 vssd1 vccd1 vccd1 _14773_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10936_ _10936_/A _10936_/B _10936_/C vssd1 vssd1 vccd1 vccd1 _10937_/C sky130_fd_sc_hd__nand3_1
XFILLER_72_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13724_ _16070_/Q _16069_/Q _16068_/Q _13723_/X vssd1 vssd1 vccd1 vccd1 _16053_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10867_ _15601_/Q _15600_/Q _15599_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _15593_/D
+ sky130_fd_sc_hd__o31a_1
X_13655_ _16043_/Q _13853_/B _13655_/C vssd1 vssd1 vccd1 vccd1 _13662_/B sky130_fd_sc_hd__and3_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12606_/A vssd1 vssd1 vccd1 vccd1 _15866_/D sky130_fd_sc_hd__clkbuf_1
X_13586_ _13580_/B _13581_/C _13583_/X _13584_/Y vssd1 vssd1 vccd1 vccd1 _13587_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _15583_/Q _10798_/B _10798_/C vssd1 vssd1 vccd1 vccd1 _10806_/B sky130_fd_sc_hd__and3_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15325_ _15337_/CLK _15325_/D vssd1 vssd1 vccd1 vccd1 _15325_/Q sky130_fd_sc_hd__dfxtp_2
X_12537_ _15856_/Q _12575_/C _12481_/X vssd1 vssd1 vccd1 vccd1 _12539_/B sky130_fd_sc_hd__a21oi_1
XFILLER_8_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15256_ _15274_/CLK _15256_/D vssd1 vssd1 vccd1 vccd1 _15256_/Q sky130_fd_sc_hd__dfxtp_1
X_12468_ _12466_/A _12466_/B _12467_/X vssd1 vssd1 vccd1 vccd1 _15843_/D sky130_fd_sc_hd__a21oi_1
XFILLER_138_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14207_ _16147_/Q _14337_/B _14207_/C vssd1 vssd1 vccd1 vccd1 _14212_/A sky130_fd_sc_hd__and3_1
X_11419_ _11417_/Y _11412_/C _11414_/X _11415_/Y vssd1 vssd1 vccd1 vccd1 _11420_/C
+ sky130_fd_sc_hd__a211o_1
X_15187_ _14408_/A _15189_/C _08335_/X vssd1 vssd1 vccd1 vccd1 _15188_/B sky130_fd_sc_hd__o21ai_1
XFILLER_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12399_ _15834_/Q _12512_/B _12399_/C vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__and3_1
XFILLER_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14138_ _16133_/Q _14137_/C _14004_/X vssd1 vssd1 vccd1 vccd1 _14139_/B sky130_fd_sc_hd__a21o_1
XFILLER_141_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14069_ _14287_/A vssd1 vssd1 vccd1 vccd1 _14069_/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_3_clk _15584_/CLK vssd1 vssd1 vccd1 vccd1 _15926_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08630_ _08630_/A vssd1 vssd1 vccd1 vccd1 _15246_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08561_ _15238_/Q _08568_/C _12609_/A vssd1 vssd1 vccd1 vccd1 _08561_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08492_ _12777_/A vssd1 vssd1 vccd1 vccd1 _10939_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09113_ _09110_/X _09111_/Y _09112_/Y _09108_/C vssd1 vssd1 vccd1 vccd1 _09115_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09044_ _09044_/A vssd1 vssd1 vccd1 vccd1 _15309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09946_ _09958_/C vssd1 vssd1 vccd1 vccd1 _09967_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _09877_/A _09877_/B vssd1 vssd1 vccd1 vccd1 _09878_/B sky130_fd_sc_hd__nor2_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08828_ _08826_/Y _08821_/C _08834_/A _08825_/Y vssd1 vssd1 vccd1 vccd1 _08834_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _15267_/Q _08769_/C _08575_/X vssd1 vssd1 vccd1 vccd1 _08759_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11778_/A _11768_/Y _11769_/Y _11765_/C vssd1 vssd1 vccd1 vccd1 _11772_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _15571_/Q _10722_/C _10663_/X vssd1 vssd1 vccd1 vccd1 _10721_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13436_/X _13438_/Y _13439_/Y _13434_/C vssd1 vssd1 vccd1 vccd1 _13442_/B
+ sky130_fd_sc_hd__o211ai_1
X_10652_ _10676_/A _10652_/B _10652_/C vssd1 vssd1 vccd1 vccd1 _10653_/A sky130_fd_sc_hd__and3_1
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13371_ _15993_/Q _13401_/C _13317_/X vssd1 vssd1 vccd1 vccd1 _13373_/B sky130_fd_sc_hd__a21oi_1
X_10583_ _10596_/C vssd1 vssd1 vccd1 vccd1 _10604_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15110_ _15110_/A _15110_/B vssd1 vssd1 vccd1 vccd1 _15111_/B sky130_fd_sc_hd__nor2_1
X_12322_ _12322_/A vssd1 vssd1 vccd1 vccd1 _15821_/D sky130_fd_sc_hd__clkbuf_1
X_16090_ _16103_/CLK _16090_/D vssd1 vssd1 vccd1 vccd1 _16090_/Q sky130_fd_sc_hd__dfxtp_2
X_15041_ _15041_/A _15041_/B vssd1 vssd1 vccd1 vccd1 _15041_/X sky130_fd_sc_hd__or2_1
X_12253_ _15811_/Q _12291_/C _12197_/X vssd1 vssd1 vccd1 vccd1 _12255_/B sky130_fd_sc_hd__a21oi_1
XFILLER_5_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ _11204_/A _11208_/C vssd1 vssd1 vccd1 vccd1 _11204_/X sky130_fd_sc_hd__or2_1
XFILLER_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ _12182_/A _12182_/B _12183_/X vssd1 vssd1 vccd1 vccd1 _15798_/D sky130_fd_sc_hd__a21oi_1
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ _11422_/A vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11066_ _15624_/Q _11121_/B _11066_/C vssd1 vssd1 vccd1 vccd1 _11066_/Y sky130_fd_sc_hd__nand3_1
X_15943_ _15196_/Q _15943_/D vssd1 vssd1 vccd1 vccd1 _15943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10017_ _15462_/Q _10024_/C _09786_/X vssd1 vssd1 vccd1 vccd1 _10017_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15874_ _07603_/A _15874_/D vssd1 vssd1 vccd1 vccd1 _15874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14825_ _14825_/A _14825_/B _14829_/A vssd1 vssd1 vccd1 vccd1 _16279_/D sky130_fd_sc_hd__nor3_1
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14756_ _16268_/Q _14755_/C _14718_/X vssd1 vssd1 vccd1 vccd1 _14757_/B sky130_fd_sc_hd__a21oi_1
X_11968_ _12000_/C vssd1 vssd1 vccd1 vccd1 _12007_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13707_ _16052_/Q _13853_/B _13707_/C vssd1 vssd1 vccd1 vccd1 _13716_/B sky130_fd_sc_hd__and3_1
X_10919_ _11783_/A vssd1 vssd1 vccd1 vccd1 _11151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11899_ _13029_/A vssd1 vssd1 vccd1 vccd1 _12129_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14687_ _14847_/A _14693_/C vssd1 vssd1 vccd1 vccd1 _14687_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13638_ _13664_/A _13638_/B _13638_/C vssd1 vssd1 vccd1 vccd1 _13639_/A sky130_fd_sc_hd__and3_1
X_16357_ _16364_/CLK _16357_/D vssd1 vssd1 vccd1 vccd1 _16357_/Q sky130_fd_sc_hd__dfxtp_1
X_13569_ _16017_/Q vssd1 vssd1 vccd1 vccd1 _13575_/C sky130_fd_sc_hd__inv_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ _15312_/CLK _15308_/D vssd1 vssd1 vccd1 vccd1 _15308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16288_ _16304_/CLK _16288_/D vssd1 vssd1 vccd1 vccd1 _16288_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_145_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15239_ _15239_/CLK _15239_/D vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfxtp_1
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09800_ _09800_/A vssd1 vssd1 vccd1 vccd1 _15426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07992_ _13937_/C _07881_/B _07991_/X vssd1 vssd1 vccd1 vccd1 _08187_/A sky130_fd_sc_hd__o21ai_2
XFILLER_101_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09731_ _09746_/A _09731_/B _09731_/C vssd1 vssd1 vccd1 vccd1 _09732_/A sky130_fd_sc_hd__and3_1
X_09662_ _15406_/Q _09700_/C _09605_/X vssd1 vssd1 vccd1 vccd1 _09664_/B sky130_fd_sc_hd__a21oi_1
XFILLER_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08613_ _13099_/A vssd1 vssd1 vccd1 vccd1 _08853_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09593_ _09825_/A vssd1 vssd1 vccd1 vccd1 _09635_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _08544_/A vssd1 vssd1 vccd1 vccd1 _15233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08475_ _08493_/C vssd1 vssd1 vccd1 vccd1 _08505_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09027_ _09061_/C vssd1 vssd1 vccd1 vccd1 _09067_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09929_ _09927_/Y _09922_/C _09934_/A _09926_/Y vssd1 vssd1 vccd1 vccd1 _09934_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12940_ _12940_/A vssd1 vssd1 vccd1 vccd1 _15919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12871_ _12906_/A _12871_/B _12871_/C vssd1 vssd1 vccd1 vccd1 _12872_/A sky130_fd_sc_hd__and3_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14610_ _14604_/Y _14605_/X _14607_/B vssd1 vssd1 vccd1 vccd1 _14611_/B sky130_fd_sc_hd__o21a_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11819_/X _11820_/Y _11821_/Y _11817_/C vssd1 vssd1 vccd1 vccd1 _11824_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15194_/Q _15590_/D vssd1 vssd1 vccd1 vccd1 _15590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11753_ _12041_/A vssd1 vssd1 vccd1 vccd1 _11986_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14541_ _14541_/A vssd1 vssd1 vccd1 vccd1 _14936_/A sky130_fd_sc_hd__buf_4
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _15568_/Q _10741_/C _10474_/X vssd1 vssd1 vccd1 vccd1 _10706_/B sky130_fd_sc_hd__a21oi_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _15722_/Q _11689_/C _11512_/X vssd1 vssd1 vccd1 vccd1 _11686_/C sky130_fd_sc_hd__a21o_1
XFILLER_81_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ _14552_/A _14472_/B _14472_/C vssd1 vssd1 vccd1 vccd1 _14473_/A sky130_fd_sc_hd__and3_1
X_16211_ _16240_/CLK _16211_/D vssd1 vssd1 vccd1 vccd1 _16211_/Q sky130_fd_sc_hd__dfxtp_1
X_10635_ _10634_/B _10634_/C _10464_/X vssd1 vssd1 vccd1 vccd1 _10636_/C sky130_fd_sc_hd__o21ai_1
X_13423_ _13679_/A vssd1 vssd1 vccd1 vccd1 _13628_/B sky130_fd_sc_hd__buf_4
XFILLER_139_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16374__23 vssd1 vssd1 vccd1 vccd1 _16374__23/HI io_oeb[6] sky130_fd_sc_hd__conb_1
XFILLER_10_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13354_ _13457_/A _13358_/C vssd1 vssd1 vccd1 vccd1 _13354_/X sky130_fd_sc_hd__or2_1
X_16142_ _16142_/CLK _16142_/D vssd1 vssd1 vccd1 vccd1 _16142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10566_ _10564_/Y _10559_/C _10572_/A _10563_/Y vssd1 vssd1 vccd1 vccd1 _10572_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12305_ _12317_/C vssd1 vssd1 vccd1 vccd1 _12326_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16073_ _16075_/CLK _16073_/D vssd1 vssd1 vccd1 vccd1 _16073_/Q sky130_fd_sc_hd__dfxtp_2
X_13285_ _15978_/Q _13291_/C _13179_/X vssd1 vssd1 vccd1 vccd1 _13285_/Y sky130_fd_sc_hd__a21oi_1
X_10497_ _15536_/Q _10609_/B _10506_/C vssd1 vssd1 vccd1 vccd1 _10497_/X sky130_fd_sc_hd__and3_1
XFILLER_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _15808_/Q _12235_/C _12063_/X vssd1 vssd1 vccd1 vccd1 _12237_/B sky130_fd_sc_hd__a21oi_1
X_15024_ _16329_/Q _15131_/B _15024_/C vssd1 vssd1 vccd1 vccd1 _15027_/B sky130_fd_sc_hd__nand3_1
XFILLER_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12167_ _15796_/Q _12223_/B _12172_/C vssd1 vssd1 vccd1 vccd1 _12167_/Y sky130_fd_sc_hd__nand3_1
XFILLER_122_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11118_ _11118_/A vssd1 vssd1 vccd1 vccd1 _15632_/D sky130_fd_sc_hd__clkbuf_1
X_12098_ _12098_/A vssd1 vssd1 vccd1 vccd1 _15785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11049_ _15622_/Q _11161_/B _11058_/C vssd1 vssd1 vccd1 vccd1 _11054_/A sky130_fd_sc_hd__and3_1
X_15926_ _15926_/CLK _15926_/D vssd1 vssd1 vccd1 vccd1 _15926_/Q sky130_fd_sc_hd__dfxtp_1
Xinput7 in1[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
XFILLER_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15857_ _07603_/A _15857_/D vssd1 vssd1 vccd1 vccd1 _15857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _15169_/A vssd1 vssd1 vccd1 vccd1 _14808_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15788_ _15195_/Q _15788_/D vssd1 vssd1 vccd1 vccd1 _15788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14739_ _14743_/C vssd1 vssd1 vccd1 vccd1 _14755_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08260_ _08260_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08260_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08191_ _08191_/A _08191_/B _08191_/C vssd1 vssd1 vccd1 vccd1 _08192_/B sky130_fd_sc_hd__nand3_1
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07975_ _07975_/A _07975_/B vssd1 vssd1 vccd1 vccd1 _07976_/B sky130_fd_sc_hd__xnor2_4
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _09727_/C vssd1 vssd1 vccd1 vccd1 _09735_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09645_ _15403_/Q _09644_/C _09467_/X vssd1 vssd1 vccd1 vccd1 _09646_/B sky130_fd_sc_hd__a21oi_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09576_ _09576_/A vssd1 vssd1 vccd1 vccd1 _15391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08535_/A _08525_/Y _08526_/Y _08519_/C vssd1 vssd1 vccd1 vccd1 _08529_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08458_ _11898_/A vssd1 vssd1 vccd1 vccd1 _14163_/A sky130_fd_sc_hd__buf_4
X_08389_ _08389_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _08404_/B sky130_fd_sc_hd__xor2_4
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10420_ _10421_/B _10421_/C _10421_/A vssd1 vssd1 vccd1 vccd1 _10422_/B sky130_fd_sc_hd__a21o_1
XFILLER_51_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10351_ _15514_/Q _10395_/C _10181_/X vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__a21oi_1
X_13070_ _13070_/A vssd1 vssd1 vccd1 vccd1 _15941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10282_ _10280_/A _10280_/B _10281_/X vssd1 vssd1 vccd1 vccd1 _15501_/D sky130_fd_sc_hd__a21oi_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12021_ _12033_/C vssd1 vssd1 vccd1 vccd1 _12042_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13972_ _13972_/A vssd1 vssd1 vccd1 vccd1 _14818_/A sky130_fd_sc_hd__buf_4
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15711_ _15794_/CLK _15711_/D vssd1 vssd1 vccd1 vccd1 _15711_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12923_ _13151_/A _12923_/B _12923_/C vssd1 vssd1 vccd1 vccd1 _12925_/B sky130_fd_sc_hd__or3_1
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15642_ _15194_/Q _15642_/D vssd1 vssd1 vccd1 vccd1 _15642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _15906_/Q _13071_/B _12854_/C vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__and3_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _12377_/A vssd1 vssd1 vccd1 vccd1 _11805_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _15655_/CLK _15573_/D vssd1 vssd1 vccd1 vccd1 _15573_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _15895_/Q _12786_/C _12668_/X vssd1 vssd1 vccd1 vccd1 _12785_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14521_/B _14520_/Y _14521_/A vssd1 vssd1 vccd1 vccd1 _14524_/Y sky130_fd_sc_hd__o21bai_1
X_11736_ _15730_/Q _11774_/C _11624_/X vssd1 vssd1 vccd1 vccd1 _11738_/B sky130_fd_sc_hd__a21oi_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14455_ _14408_/X _14453_/B _14454_/Y vssd1 vssd1 vccd1 vccd1 _16194_/D sky130_fd_sc_hd__o21a_1
X_11667_ _11780_/A _11670_/C vssd1 vssd1 vccd1 vccd1 _11667_/X sky130_fd_sc_hd__or2_1
X_13406_ _13457_/A _13408_/C vssd1 vssd1 vccd1 vccd1 _13406_/X sky130_fd_sc_hd__or2_1
X_10618_ _15555_/Q _10623_/C _10562_/X vssd1 vssd1 vccd1 vccd1 _10618_/Y sky130_fd_sc_hd__a21oi_1
X_14386_ _14386_/A _14386_/B _14386_/C vssd1 vssd1 vccd1 vccd1 _14387_/C sky130_fd_sc_hd__nand3_1
X_11598_ _11598_/A vssd1 vssd1 vccd1 vccd1 _15706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16125_ _16143_/CLK _16125_/D vssd1 vssd1 vccd1 vccd1 _16125_/Q sky130_fd_sc_hd__dfxtp_1
X_10549_ _15543_/Q _10778_/B _10549_/C vssd1 vssd1 vccd1 vccd1 _10549_/Y sky130_fd_sc_hd__nand3_1
X_13337_ _13333_/X _13334_/Y _13336_/Y _13331_/C vssd1 vssd1 vccd1 vccd1 _13339_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_128_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16056_ _16075_/CLK _16056_/D vssd1 vssd1 vccd1 vccd1 _16056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13268_ _15976_/Q _13374_/B _13276_/C vssd1 vssd1 vccd1 vccd1 _13272_/B sky130_fd_sc_hd__nand3_1
XFILLER_142_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15007_ _15086_/A vssd1 vssd1 vccd1 vccd1 _15007_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12219_ _12226_/A _12219_/B _12219_/C vssd1 vssd1 vccd1 vccd1 _12220_/A sky130_fd_sc_hd__and3_1
X_13199_ _13199_/A _13202_/C vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__or2_1
XFILLER_97_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07760_ _15926_/Q vssd1 vssd1 vccd1 vccd1 _12983_/A sky130_fd_sc_hd__clkinv_2
Xclkbuf_1_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15909_ _15196_/Q _15909_/D vssd1 vssd1 vccd1 vccd1 _15909_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07691_ _07688_/X _07698_/C _07690_/X vssd1 vssd1 vccd1 vccd1 _07692_/B sky130_fd_sc_hd__o21ai_1
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09430_ _15370_/Q _09663_/B _09438_/C vssd1 vssd1 vccd1 vccd1 _09435_/A sky130_fd_sc_hd__and3_1
XFILLER_65_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _09536_/A vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08312_ _08312_/A _08312_/B vssd1 vssd1 vccd1 vccd1 _08312_/Y sky130_fd_sc_hd__nor2_1
X_09292_ _13598_/A vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__buf_2
XANTENNA_12 _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08243_/A vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__inv_2
XANTENNA_23 _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 hold25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ _08174_/A _08159_/A vssd1 vssd1 vccd1 vccd1 _08270_/B sky130_fd_sc_hd__or2b_1
XFILLER_119_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07958_ _07920_/A _07920_/B _07957_/Y vssd1 vssd1 vccd1 vccd1 _07977_/A sky130_fd_sc_hd__o21ai_4
XFILLER_101_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07889_ _15422_/Q _07890_/B vssd1 vssd1 vccd1 vccd1 _07891_/A sky130_fd_sc_hd__or2_1
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09628_ _15401_/Q _09740_/B _09638_/C vssd1 vssd1 vccd1 vccd1 _09628_/X sky130_fd_sc_hd__and3_1
XFILLER_55_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09559_ _09557_/X _09558_/Y _09553_/B _09554_/C vssd1 vssd1 vccd1 vccd1 _09561_/B
+ sky130_fd_sc_hd__o211ai_1
X_12570_ _15861_/Q _12575_/C _12569_/X vssd1 vssd1 vccd1 vccd1 _12570_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11521_ _11518_/X _11520_/Y _11515_/B _11516_/C vssd1 vssd1 vccd1 vccd1 _11523_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11452_ _15686_/Q _11457_/C _11222_/X vssd1 vssd1 vccd1 vccd1 _11454_/C sky130_fd_sc_hd__a21o_1
X_14240_ _14459_/A vssd1 vssd1 vccd1 vccd1 _14240_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10403_ _10401_/A _10401_/B _10402_/X vssd1 vssd1 vccd1 vccd1 _15519_/D sky130_fd_sc_hd__a21oi_1
X_14171_ _16140_/Q _14256_/B _14171_/C vssd1 vssd1 vccd1 vccd1 _14179_/A sky130_fd_sc_hd__and3_1
X_11383_ _11382_/B _11382_/C _11327_/X vssd1 vssd1 vccd1 vccd1 _11384_/C sky130_fd_sc_hd__o21ai_1
XFILLER_124_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10334_ _15511_/Q _10331_/C _10333_/X vssd1 vssd1 vccd1 vccd1 _10335_/B sky130_fd_sc_hd__a21oi_1
X_13122_ _15950_/Q _13286_/B _13127_/C vssd1 vssd1 vccd1 vccd1 _13122_/Y sky130_fd_sc_hd__nand3_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13053_ _13051_/X _13052_/Y _13048_/B _13049_/C vssd1 vssd1 vccd1 vccd1 _13055_/B
+ sky130_fd_sc_hd__o211ai_1
X_10265_ _10263_/Y _10259_/C _10261_/X _10262_/Y vssd1 vssd1 vccd1 vccd1 _10266_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ _12010_/A _12002_/Y _12003_/Y _11997_/C vssd1 vssd1 vccd1 vccd1 _12006_/B
+ sky130_fd_sc_hd__o211a_1
X_10196_ _10196_/A vssd1 vssd1 vccd1 vccd1 _15488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13955_ _13953_/A _13953_/B _13952_/Y _13954_/Y vssd1 vssd1 vccd1 vccd1 _16093_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12906_ _12906_/A _12906_/B _12906_/C vssd1 vssd1 vccd1 vccd1 _12907_/A sky130_fd_sc_hd__and3_1
XFILLER_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _16086_/Q _13885_/C _14088_/B vssd1 vssd1 vccd1 vccd1 _13886_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15625_ _15194_/Q _15625_/D vssd1 vssd1 vccd1 vccd1 _15625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12837_/A vssd1 vssd1 vccd1 vccd1 _15902_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _15655_/CLK _15556_/D vssd1 vssd1 vccd1 vccd1 _15556_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _15892_/Q _12805_/C _12767_/X vssd1 vssd1 vccd1 vccd1 _12770_/B sky130_fd_sc_hd__a21oi_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _16211_/Q _14587_/B _14513_/C vssd1 vssd1 vccd1 vccd1 _14510_/B sky130_fd_sc_hd__nand3_1
X_11719_ _15727_/Q _11719_/B _11719_/C vssd1 vssd1 vccd1 vccd1 _11727_/B sky130_fd_sc_hd__and3_1
X_15487_ _15224_/Q _15487_/D vssd1 vssd1 vccd1 vccd1 _15487_/Q sky130_fd_sc_hd__dfxtp_1
X_12699_ _12869_/A _12699_/B _12699_/C vssd1 vssd1 vccd1 vccd1 _12701_/B sky130_fd_sc_hd__or3_1
XFILLER_30_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14438_ _14431_/B _14432_/C _14442_/A _14436_/Y vssd1 vssd1 vccd1 vccd1 _14442_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_143_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14369_ _14368_/X _14366_/B _14316_/X vssd1 vssd1 vccd1 vccd1 _14369_/Y sky130_fd_sc_hd__a21oi_1
X_16108_ _16119_/CLK _16108_/D vssd1 vssd1 vccd1 vccd1 _16108_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16039_ _16040_/CLK _16039_/D vssd1 vssd1 vccd1 vccd1 _16039_/Q sky130_fd_sc_hd__dfxtp_1
X_08930_ _15293_/Q _08931_/C _08929_/X vssd1 vssd1 vccd1 vccd1 _08930_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08861_ _08859_/X _08860_/Y _08856_/B _08857_/C vssd1 vssd1 vccd1 vccd1 _08863_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_111_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07812_ _14466_/C _08059_/B vssd1 vssd1 vccd1 vccd1 _07818_/A sky130_fd_sc_hd__xnor2_1
XFILLER_97_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08792_ _08823_/C vssd1 vssd1 vccd1 vccd1 _08831_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_85_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07743_ _16296_/Q vssd1 vssd1 vccd1 vccd1 _08106_/A sky130_fd_sc_hd__inv_2
XFILLER_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07674_ _07674_/A vssd1 vssd1 vccd1 vccd1 _15001_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09413_ _09419_/B _09413_/B vssd1 vssd1 vccd1 vccd1 _09415_/A sky130_fd_sc_hd__or2_1
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09344_ _09342_/Y _09337_/C _09339_/X _09340_/Y vssd1 vssd1 vccd1 vccd1 _09345_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ _09275_/A vssd1 vssd1 vccd1 vccd1 _15345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08226_ _08226_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _08305_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _08966_/A _07937_/B _08156_/Y vssd1 vssd1 vccd1 vccd1 _08173_/B sky130_fd_sc_hd__o21a_1
XFILLER_107_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08088_ _15575_/Q _08088_/B vssd1 vssd1 vccd1 vccd1 _08088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10050_ _10048_/A _10048_/B _10049_/X vssd1 vssd1 vccd1 vccd1 _15465_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13740_ _13738_/X _13739_/Y _13734_/B _13735_/C vssd1 vssd1 vccd1 vccd1 _13742_/B
+ sky130_fd_sc_hd__o211ai_1
X_10952_ _10950_/Y _10944_/C _10946_/X _10949_/Y vssd1 vssd1 vccd1 vccd1 _10953_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ _13675_/C vssd1 vssd1 vccd1 vccd1 _13686_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10883_ _15597_/Q _10890_/C _10655_/X vssd1 vssd1 vccd1 vccd1 _10883_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15410_ _15483_/CLK _15410_/D vssd1 vssd1 vccd1 vccd1 _15410_/Q sky130_fd_sc_hd__dfxtp_1
X_12622_ _12622_/A vssd1 vssd1 vccd1 vccd1 _15868_/D sky130_fd_sc_hd__clkbuf_1
X_15341_ _15368_/CLK _15341_/D vssd1 vssd1 vccd1 vccd1 _15341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12553_ _15859_/Q _12554_/C _12384_/X vssd1 vssd1 vccd1 vccd1 _12553_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11504_ _11528_/C vssd1 vssd1 vccd1 vccd1 _11541_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15272_ _15282_/CLK _15272_/D vssd1 vssd1 vccd1 vccd1 _15272_/Q sky130_fd_sc_hd__dfxtp_1
X_12484_ _12518_/A _12484_/B _12488_/A vssd1 vssd1 vccd1 vccd1 _15846_/D sky130_fd_sc_hd__nor3_1
XFILLER_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14223_ _14223_/A _14223_/B vssd1 vssd1 vccd1 vccd1 _14223_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11435_ _11435_/A _11435_/B vssd1 vssd1 vccd1 vccd1 _11439_/C sky130_fd_sc_hd__nor2_1
X_11366_ _11366_/A vssd1 vssd1 vccd1 vccd1 _15670_/D sky130_fd_sc_hd__clkbuf_1
X_14154_ _14061_/X _14153_/X _14146_/B _13969_/X vssd1 vssd1 vccd1 vccd1 _14155_/B
+ sky130_fd_sc_hd__a31o_1
X_10317_ _15509_/Q _10317_/B _10325_/C vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__and3_1
X_13105_ _13105_/A _13105_/B _13105_/C vssd1 vssd1 vccd1 vccd1 _13106_/C sky130_fd_sc_hd__nand3_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11297_ _15661_/Q _11298_/C _11237_/X vssd1 vssd1 vccd1 vccd1 _11297_/Y sky130_fd_sc_hd__a21oi_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _14085_/A vssd1 vssd1 vccd1 vccd1 _16119_/D sky130_fd_sc_hd__clkbuf_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _15498_/Q _10256_/C _10075_/X vssd1 vssd1 vccd1 vccd1 _10248_/Y sky130_fd_sc_hd__a21oi_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _15951_/Q _15953_/Q _15952_/Q _12981_/X vssd1 vssd1 vccd1 vccd1 _15936_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_78_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10179_ _10199_/C vssd1 vssd1 vccd1 vccd1 _10214_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14987_ hold5/A _15031_/B _14994_/C vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__and3_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13938_ _13980_/A _13938_/B _13942_/A vssd1 vssd1 vccd1 vccd1 _16090_/D sky130_fd_sc_hd__nor3_1
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13869_ _16215_/Q vssd1 vssd1 vccd1 vccd1 _13874_/C sky130_fd_sc_hd__inv_2
X_15608_ _15194_/Q _15608_/D vssd1 vssd1 vccd1 vccd1 _15608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15539_ _15539_/CLK _15539_/D vssd1 vssd1 vccd1 vccd1 _15539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ _09924_/A vssd1 vssd1 vccd1 vccd1 _09290_/B sky130_fd_sc_hd__buf_2
X_08011_ _08207_/A _08011_/B vssd1 vssd1 vccd1 vccd1 _08014_/A sky130_fd_sc_hd__or2_1
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09962_ _09977_/A _09962_/B _09962_/C vssd1 vssd1 vccd1 vccd1 _09963_/A sky130_fd_sc_hd__and3_1
XFILLER_116_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08913_ _09778_/A vssd1 vssd1 vccd1 vccd1 _08913_/X sky130_fd_sc_hd__clkbuf_2
X_09893_ _10181_/A vssd1 vssd1 vccd1 vccd1 _09893_/X sky130_fd_sc_hd__clkbuf_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08844_ _15270_/Q vssd1 vssd1 vccd1 vccd1 _08859_/C sky130_fd_sc_hd__inv_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08775_ _15269_/Q _08775_/B _08775_/C vssd1 vssd1 vccd1 vccd1 _08783_/B sky130_fd_sc_hd__and3_1
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07726_ _15279_/Q _15261_/Q vssd1 vssd1 vccd1 vccd1 _07727_/B sky130_fd_sc_hd__or2_1
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07657_ _14993_/A vssd1 vssd1 vccd1 vccd1 _14755_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09327_ _15355_/Q _09334_/C _09212_/X vssd1 vssd1 vccd1 vccd1 _09327_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09258_ _09278_/C vssd1 vssd1 vccd1 vccd1 _09290_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08209_ _08209_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08219_/A sky130_fd_sc_hd__xor2_4
X_09189_ _10341_/A vssd1 vssd1 vccd1 vccd1 _09419_/A sky130_fd_sc_hd__clkbuf_2
X_11220_ _11220_/A _11220_/B _11225_/A vssd1 vssd1 vccd1 vccd1 _15648_/D sky130_fd_sc_hd__nor3_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11151_ _11151_/A _11151_/B _11151_/C vssd1 vssd1 vccd1 vccd1 _11153_/B sky130_fd_sc_hd__or3_1
XFILLER_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10102_ _15473_/Q _10102_/B _10106_/C vssd1 vssd1 vccd1 vccd1 _10102_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _15626_/Q _11313_/B _11086_/C vssd1 vssd1 vccd1 vccd1 _11082_/Y sky130_fd_sc_hd__nand3_1
XFILLER_95_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10033_ _10029_/X _10031_/Y _10032_/Y _10027_/C vssd1 vssd1 vccd1 vccd1 _10035_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14910_ _14910_/A vssd1 vssd1 vccd1 vccd1 _16298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15890_ _15890_/CLK _15890_/D vssd1 vssd1 vccd1 vccd1 _15890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14841_ _14841_/A _14841_/B vssd1 vssd1 vccd1 vccd1 _14842_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14772_ _14970_/A vssd1 vssd1 vccd1 vccd1 _14772_/X sky130_fd_sc_hd__clkbuf_2
X_11984_ _15769_/Q _12099_/B _11986_/C vssd1 vssd1 vccd1 vccd1 _11984_/X sky130_fd_sc_hd__and3_1
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13723_ _13723_/A vssd1 vssd1 vccd1 vccd1 _13723_/X sky130_fd_sc_hd__buf_2
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10935_ _10936_/B _10936_/C _10936_/A vssd1 vssd1 vccd1 vccd1 _10937_/B sky130_fd_sc_hd__a21o_1
XFILLER_72_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13654_ _13654_/A vssd1 vssd1 vccd1 vccd1 _13853_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10866_ _10866_/A vssd1 vssd1 vccd1 vccd1 _15592_/D sky130_fd_sc_hd__clkbuf_1
X_12605_ _12621_/A _12605_/B _12605_/C vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__and3_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13583_/X _13584_/Y _13580_/B _13581_/C vssd1 vssd1 vccd1 vccd1 _13587_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_129_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ _10797_/A _10797_/B _10801_/B vssd1 vssd1 vccd1 vccd1 _15581_/D sky130_fd_sc_hd__nor3_1
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _15368_/CLK _15324_/D vssd1 vssd1 vccd1 vccd1 _15324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12536_ _12568_/C vssd1 vssd1 vccd1 vccd1 _12575_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15255_ _15274_/CLK _15255_/D vssd1 vssd1 vccd1 vccd1 _15255_/Q sky130_fd_sc_hd__dfxtp_1
X_12467_ _12636_/A _12471_/C vssd1 vssd1 vccd1 vccd1 _12467_/X sky130_fd_sc_hd__or2_1
X_14206_ _16147_/Q _14228_/C _14069_/X vssd1 vssd1 vccd1 vccd1 _14208_/B sky130_fd_sc_hd__a21oi_1
X_11418_ _11414_/X _11415_/Y _11417_/Y _11412_/C vssd1 vssd1 vccd1 vccd1 _11420_/B
+ sky130_fd_sc_hd__o211ai_1
X_15186_ _15186_/A _15189_/C vssd1 vssd1 vccd1 vccd1 _15188_/A sky130_fd_sc_hd__and2_1
X_12398_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__buf_2
XFILLER_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ _16133_/Q _14137_/B _14137_/C vssd1 vssd1 vccd1 vccd1 _14137_/X sky130_fd_sc_hd__and3_1
X_11349_ _11347_/X _11348_/Y _11343_/B _11344_/C vssd1 vssd1 vccd1 vccd1 _11351_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_99_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14068_ _14093_/C vssd1 vssd1 vccd1 vccd1 _14099_/C sky130_fd_sc_hd__clkbuf_2
X_13019_ _13025_/A _13017_/Y _13018_/Y _13014_/C vssd1 vssd1 vccd1 vccd1 _13021_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08560_ _15238_/Q _10939_/C _08560_/C vssd1 vssd1 vccd1 vccd1 _08560_/X sky130_fd_sc_hd__and3_1
X_08491_ input3/X vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__buf_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09112_ _15320_/Q _09285_/B _09117_/C vssd1 vssd1 vccd1 vccd1 _09112_/Y sky130_fd_sc_hd__nand3_1
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09043_ _09058_/A _09043_/B _09043_/C vssd1 vssd1 vccd1 vccd1 _09044_/A sky130_fd_sc_hd__and3_1
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ _15449_/Q vssd1 vssd1 vccd1 vccd1 _09958_/C sky130_fd_sc_hd__inv_2
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09883_/B _09876_/B vssd1 vssd1 vccd1 vccd1 _09878_/A sky130_fd_sc_hd__or2_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08827_ _08834_/A _08825_/Y _08826_/Y _08821_/C vssd1 vssd1 vccd1 vccd1 _08829_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _15267_/Q _08872_/B _08769_/C vssd1 vssd1 vccd1 vccd1 _08758_/X sky130_fd_sc_hd__and3_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _12758_/A vssd1 vssd1 vccd1 vccd1 _14970_/A sky130_fd_sc_hd__buf_4
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08682_/B _08683_/C _08686_/X _08687_/Y vssd1 vssd1 vccd1 vccd1 _08690_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _15571_/Q _10888_/B _10722_/C vssd1 vssd1 vccd1 vccd1 _10720_/X sky130_fd_sc_hd__and3_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10651_ _10651_/A _10651_/B _10651_/C vssd1 vssd1 vccd1 vccd1 _10652_/C sky130_fd_sc_hd__nand3_1
XFILLER_139_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10582_ _15548_/Q vssd1 vssd1 vccd1 vccd1 _10596_/C sky130_fd_sc_hd__inv_2
X_13370_ _13394_/C vssd1 vssd1 vccd1 vccd1 _13401_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_139_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12321_ _12337_/A _12321_/B _12321_/C vssd1 vssd1 vccd1 vccd1 _12322_/A sky130_fd_sc_hd__and3_1
XFILLER_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15040_ _15040_/A _15040_/B vssd1 vssd1 vccd1 vccd1 _15041_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12252_ _12284_/C vssd1 vssd1 vccd1 vccd1 _12291_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_135_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11203_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _11208_/C sky130_fd_sc_hd__nor2_1
X_12183_ _12352_/A _12187_/C vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__or2_1
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11134_ _11134_/A vssd1 vssd1 vccd1 vccd1 _15634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11065_ _15625_/Q _11066_/C _10948_/X vssd1 vssd1 vccd1 vccd1 _11065_/Y sky130_fd_sc_hd__a21oi_1
X_15942_ _15196_/Q _15942_/D vssd1 vssd1 vccd1 vccd1 _15942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10016_ _15462_/Q _10074_/B _10016_/C vssd1 vssd1 vccd1 vccd1 _10016_/X sky130_fd_sc_hd__and3_1
XFILLER_95_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15873_ _07603_/A _15873_/D vssd1 vssd1 vccd1 vccd1 _15873_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14824_ _16283_/Q _14977_/B _14826_/C vssd1 vssd1 vccd1 vccd1 _14829_/A sky130_fd_sc_hd__and3_1
X_14755_ _16268_/Q _14755_/B _14755_/C vssd1 vssd1 vccd1 vccd1 _14757_/A sky130_fd_sc_hd__and3_1
X_11967_ _11986_/C vssd1 vssd1 vccd1 vccd1 _12000_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13706_ _13730_/A _13706_/B _13711_/B vssd1 vssd1 vccd1 vccd1 _16049_/D sky130_fd_sc_hd__nor3_1
X_10918_ _10978_/A vssd1 vssd1 vccd1 vccd1 _10960_/A sky130_fd_sc_hd__clkbuf_2
X_14686_ _14679_/A _14683_/B _14646_/X vssd1 vssd1 vccd1 vccd1 _14693_/C sky130_fd_sc_hd__o21a_1
X_11898_ _11898_/A vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__buf_2
XFILLER_60_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13637_ _13631_/B _13632_/C _13634_/X _13635_/Y vssd1 vssd1 vccd1 vccd1 _13638_/C
+ sky130_fd_sc_hd__a211o_1
X_10849_ _15591_/Q _10855_/C _10848_/X vssd1 vssd1 vccd1 vccd1 _10849_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16356_ _16364_/CLK _16356_/D vssd1 vssd1 vccd1 vccd1 _16356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ _16043_/Q _16042_/Q _16041_/Q _13467_/X vssd1 vssd1 vccd1 vccd1 _16026_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15307_ _16327_/CLK _15307_/D vssd1 vssd1 vccd1 vccd1 _15307_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_145_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12519_ _15853_/Q _12575_/B _12519_/C vssd1 vssd1 vccd1 vccd1 _12527_/B sky130_fd_sc_hd__and3_1
X_16287_ _16304_/CLK _16287_/D vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfxtp_1
X_13499_ _16015_/Q _13504_/C _13342_/X vssd1 vssd1 vccd1 vccd1 _13499_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15238_ _15239_/CLK _15238_/D vssd1 vssd1 vccd1 vccd1 _15238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _15169_/A _15169_/B _15169_/C vssd1 vssd1 vccd1 vccd1 _15170_/A sky130_fd_sc_hd__and3_1
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07991_ _07991_/A _07991_/B vssd1 vssd1 vccd1 vccd1 _07991_/X sky130_fd_sc_hd__or2_1
XFILLER_140_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09730_ _09724_/B _09725_/C _09727_/X _09728_/Y vssd1 vssd1 vccd1 vccd1 _09731_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_101_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09661_ _09692_/C vssd1 vssd1 vccd1 vccd1 _09700_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_95_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08612_ _10354_/A vssd1 vssd1 vccd1 vccd1 _13099_/A sky130_fd_sc_hd__buf_4
X_09592_ _10169_/A vssd1 vssd1 vccd1 vccd1 _09825_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08543_ _08580_/A _08543_/B _08543_/C vssd1 vssd1 vccd1 vccd1 _08544_/A sky130_fd_sc_hd__and3_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08474_ _15351_/Q vssd1 vssd1 vccd1 vccd1 _08493_/C sky130_fd_sc_hd__inv_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09026_ _09047_/C vssd1 vssd1 vccd1 vccd1 _09061_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09928_ _09934_/A _09926_/Y _09927_/Y _09922_/C vssd1 vssd1 vccd1 vccd1 _09930_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09859_ _09859_/A vssd1 vssd1 vccd1 vccd1 _15435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12870_ _12869_/B _12869_/C _12758_/X vssd1 vssd1 vccd1 vccd1 _12871_/C sky130_fd_sc_hd__o21ai_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11821_ _15742_/Q _11938_/B _11827_/C vssd1 vssd1 vccd1 vccd1 _11821_/Y sky130_fd_sc_hd__nand3_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _16088_/Q _16087_/Q _16086_/Q _14421_/X vssd1 vssd1 vccd1 vccd1 _16215_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _15733_/Q _11754_/C _11526_/X vssd1 vssd1 vccd1 vccd1 _11752_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10734_/C vssd1 vssd1 vccd1 vccd1 _10741_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14471_/A _14471_/B _14471_/C vssd1 vssd1 vccd1 vccd1 _14472_/C sky130_fd_sc_hd__nand3_1
X_11683_ _15722_/Q _11797_/B _11689_/C vssd1 vssd1 vccd1 vccd1 _11686_/B sky130_fd_sc_hd__nand3_1
XFILLER_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16240_/CLK _16210_/D vssd1 vssd1 vccd1 vccd1 _16210_/Q sky130_fd_sc_hd__dfxtp_1
X_13422_ _13612_/A vssd1 vssd1 vccd1 vccd1 _13481_/A sky130_fd_sc_hd__clkbuf_2
X_10634_ _10863_/A _10634_/B _10634_/C vssd1 vssd1 vccd1 vccd1 _10636_/B sky130_fd_sc_hd__or3_1
XFILLER_10_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _16142_/CLK _16141_/D vssd1 vssd1 vccd1 vccd1 _16141_/Q sky130_fd_sc_hd__dfxtp_1
X_13353_ _13353_/A _13353_/B vssd1 vssd1 vccd1 vccd1 _13358_/C sky130_fd_sc_hd__nor2_1
X_10565_ _10572_/A _10563_/Y _10564_/Y _10559_/C vssd1 vssd1 vccd1 vccd1 _10567_/B
+ sky130_fd_sc_hd__o211a_1
X_12304_ _12304_/A vssd1 vssd1 vccd1 vccd1 _12317_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16072_ _16129_/CLK _16072_/D vssd1 vssd1 vccd1 vccd1 _16072_/Q sky130_fd_sc_hd__dfxtp_2
X_13284_ _15978_/Q _13333_/B _13291_/C vssd1 vssd1 vccd1 vccd1 _13284_/X sky130_fd_sc_hd__and3_1
XFILLER_5_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10496_ _10496_/A vssd1 vssd1 vccd1 vccd1 _15534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15023_ _15023_/A _15023_/B _15027_/A vssd1 vssd1 vccd1 vccd1 _16324_/D sky130_fd_sc_hd__nor3_1
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12235_ _15808_/Q _12291_/B _12235_/C vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__and3_1
XFILLER_135_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12166_ _15797_/Q _12172_/C _12048_/X vssd1 vssd1 vccd1 vccd1 _12166_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11117_ _11133_/A _11117_/B _11117_/C vssd1 vssd1 vccd1 vccd1 _11118_/A sky130_fd_sc_hd__and3_1
XFILLER_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12097_ _12112_/A _12097_/B _12097_/C vssd1 vssd1 vccd1 vccd1 _12098_/A sky130_fd_sc_hd__and3_1
X_11048_ _15622_/Q _11086_/C _11047_/X vssd1 vssd1 vccd1 vccd1 _11050_/B sky130_fd_sc_hd__a21oi_1
X_15925_ _07603_/A _15925_/D vssd1 vssd1 vccd1 vccd1 _15925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 in1[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_8
X_15856_ _07603_/A _15856_/D vssd1 vssd1 vccd1 vccd1 _15856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14807_ _14963_/A _14811_/C vssd1 vssd1 vccd1 vccd1 _14810_/A sky130_fd_sc_hd__and2_1
XFILLER_92_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15787_ _15195_/Q _15787_/D vssd1 vssd1 vccd1 vccd1 _15787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12999_ _12993_/B _12994_/C _12996_/X _12997_/Y vssd1 vssd1 vccd1 vccd1 _13000_/C
+ sky130_fd_sc_hd__a211o_1
X_14738_ _16251_/Q vssd1 vssd1 vccd1 vccd1 _14743_/C sky130_fd_sc_hd__inv_2
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14669_ _14748_/A _14669_/B _14669_/C vssd1 vssd1 vccd1 vccd1 _14670_/A sky130_fd_sc_hd__and3_1
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08190_ _08191_/A _08191_/B _08191_/C vssd1 vssd1 vccd1 vccd1 _08295_/A sky130_fd_sc_hd__a21o_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16339_ _16359_/CLK _16339_/D vssd1 vssd1 vccd1 vccd1 _16339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07974_ _07974_/A _07974_/B vssd1 vssd1 vccd1 vccd1 _07975_/B sky130_fd_sc_hd__nor2_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09713_ _15413_/Q vssd1 vssd1 vccd1 vccd1 _09727_/C sky130_fd_sc_hd__inv_2
XFILLER_68_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09644_ _15403_/Q _09644_/B _09644_/C vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__and3_1
XFILLER_83_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ _09575_/A _09575_/B _09575_/C vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__and3_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _15231_/Q _10965_/C _08532_/C vssd1 vssd1 vccd1 vccd1 _08526_/Y sky130_fd_sc_hd__nand3_1
XFILLER_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08457_ _08457_/A vssd1 vssd1 vccd1 vccd1 _15220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _08388_/A _08388_/B vssd1 vssd1 vccd1 vccd1 _08389_/B sky130_fd_sc_hd__xor2_4
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _10389_/C vssd1 vssd1 vccd1 vccd1 _10395_/C sky130_fd_sc_hd__clkbuf_2
X_09009_ hold29/A _09008_/C _08888_/X vssd1 vssd1 vccd1 vccd1 _09010_/B sky130_fd_sc_hd__a21oi_1
XFILLER_124_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10281_ _10338_/A _10284_/C vssd1 vssd1 vccd1 vccd1 _10281_/X sky130_fd_sc_hd__or2_1
XFILLER_105_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ _15773_/Q vssd1 vssd1 vccd1 vccd1 _12033_/C sky130_fd_sc_hd__inv_2
XFILLER_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13971_ _13971_/A _13971_/B vssd1 vssd1 vccd1 vccd1 _16097_/D sky130_fd_sc_hd__nor2_1
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15710_ _15728_/CLK _15710_/D vssd1 vssd1 vccd1 vccd1 _15710_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12922_ input8/X vssd1 vssd1 vccd1 vccd1 _13151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15641_ _15194_/Q _15641_/D vssd1 vssd1 vccd1 vccd1 _15641_/Q sky130_fd_sc_hd__dfxtp_1
X_12853_ _12853_/A vssd1 vssd1 vccd1 vccd1 _13071_/B sky130_fd_sc_hd__buf_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11804_ _15741_/Q _11863_/B _11804_/C vssd1 vssd1 vccd1 vccd1 _11804_/X sky130_fd_sc_hd__and3_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15655_/CLK _15572_/D vssd1 vssd1 vccd1 vccd1 _15572_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _15895_/Q _12947_/B _12786_/C vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__and3_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14521_/A _14521_/B _14520_/Y _14522_/Y vssd1 vssd1 vccd1 vccd1 _16210_/D
+ sky130_fd_sc_hd__o31a_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11735_ _11767_/C vssd1 vssd1 vccd1 vccd1 _11774_/C sky130_fd_sc_hd__clkbuf_2
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _14533_/A _14454_/B vssd1 vssd1 vccd1 vccd1 _14454_/Y sky130_fd_sc_hd__nor2_1
X_11666_ _11666_/A _11666_/B vssd1 vssd1 vccd1 vccd1 _11670_/C sky130_fd_sc_hd__nor2_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13405_ _13405_/A _13405_/B vssd1 vssd1 vccd1 vccd1 _13408_/C sky130_fd_sc_hd__nor2_1
X_10617_ _15555_/Q _10734_/B _10617_/C vssd1 vssd1 vccd1 vccd1 _10627_/A sky130_fd_sc_hd__and3_1
X_14385_ _14386_/B _14386_/C _14386_/A vssd1 vssd1 vccd1 vccd1 _14387_/B sky130_fd_sc_hd__a21o_1
X_11597_ _11597_/A _11597_/B _11597_/C vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__and3_1
X_16124_ _16124_/CLK _16124_/D vssd1 vssd1 vccd1 vccd1 _16124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13336_ _15986_/Q _13543_/B _13341_/C vssd1 vssd1 vccd1 vccd1 _13336_/Y sky130_fd_sc_hd__nand3_1
X_10548_ _10548_/A vssd1 vssd1 vccd1 vccd1 _10778_/B sky130_fd_sc_hd__buf_2
XFILLER_127_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16055_ _16075_/CLK _16055_/D vssd1 vssd1 vccd1 vccd1 _16055_/Q sky130_fd_sc_hd__dfxtp_2
X_13267_ _13348_/A _13267_/B _13272_/A vssd1 vssd1 vccd1 vccd1 _15973_/D sky130_fd_sc_hd__nor3_1
X_10479_ _15533_/Q _10484_/C _10357_/X vssd1 vssd1 vccd1 vccd1 _10481_/C sky130_fd_sc_hd__a21o_1
X_15006_ _15152_/A _15010_/C vssd1 vssd1 vccd1 vccd1 _15009_/A sky130_fd_sc_hd__and2_1
X_12218_ _12216_/Y _12212_/C _12214_/X _12215_/Y vssd1 vssd1 vccd1 vccd1 _12219_/C
+ sky130_fd_sc_hd__a211o_1
X_13198_ _13198_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13202_/C sky130_fd_sc_hd__nor2_1
X_12149_ _12149_/A vssd1 vssd1 vccd1 vccd1 _15793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15908_ _15926_/CLK _15908_/D vssd1 vssd1 vccd1 vccd1 _15908_/Q sky130_fd_sc_hd__dfxtp_1
X_07690_ _15169_/A vssd1 vssd1 vccd1 vccd1 _07690_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15839_ _15907_/CLK _15839_/D vssd1 vssd1 vccd1 vccd1 _15839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09360_ _09358_/A _09358_/B _09359_/X vssd1 vssd1 vccd1 vccd1 _15358_/D sky130_fd_sc_hd__a21oi_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08311_ _08311_/A _08311_/B vssd1 vssd1 vccd1 vccd1 _08315_/A sky130_fd_sc_hd__xnor2_1
X_09291_ _15349_/Q _09297_/C _09118_/X vssd1 vssd1 vccd1 vccd1 _09291_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _08242_/A _08242_/B vssd1 vssd1 vccd1 vccd1 _08246_/A sky130_fd_sc_hd__and2_1
XFILLER_138_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_24 _14466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _13720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08173_ _08173_/A _08173_/B vssd1 vssd1 vccd1 vccd1 _08270_/A sky130_fd_sc_hd__or2_1
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07957_ _15764_/Q _07957_/B vssd1 vssd1 vccd1 vccd1 _07957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07888_ _07986_/A _07888_/B vssd1 vssd1 vccd1 vccd1 _07890_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _09627_/A vssd1 vssd1 vccd1 vccd1 _15399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09558_ _15390_/Q _09565_/C _09497_/X vssd1 vssd1 vccd1 vccd1 _09558_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08509_ _08509_/A vssd1 vssd1 vccd1 vccd1 _15229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09489_ _15380_/Q _09721_/B _09496_/C vssd1 vssd1 vccd1 vccd1 _09493_/B sky130_fd_sc_hd__nand3_1
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11520_ _15696_/Q _11528_/C _11519_/X vssd1 vssd1 vccd1 vccd1 _11520_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ _15686_/Q _11510_/B _11457_/C vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__nand3_1
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10402_ _10629_/A _10405_/C vssd1 vssd1 vccd1 vccd1 _10402_/X sky130_fd_sc_hd__or2_1
X_14170_ _14170_/A vssd1 vssd1 vccd1 vccd1 _16136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11382_ _11439_/A _11382_/B _11382_/C vssd1 vssd1 vccd1 vccd1 _11384_/B sky130_fd_sc_hd__or3_1
X_13121_ _14593_/B vssd1 vssd1 vccd1 vccd1 _13286_/B sky130_fd_sc_hd__clkbuf_4
X_10333_ _11488_/A vssd1 vssd1 vccd1 vccd1 _10333_/X sky130_fd_sc_hd__buf_2
XFILLER_124_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ _15940_/Q _13059_/C _13275_/A vssd1 vssd1 vccd1 vccd1 _13052_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10264_ _10261_/X _10262_/Y _10263_/Y _10259_/C vssd1 vssd1 vccd1 vccd1 _10266_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_127_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12003_ _15770_/Q _12174_/B _12007_/C vssd1 vssd1 vccd1 vccd1 _12003_/Y sky130_fd_sc_hd__nand3_1
X_10195_ _10210_/A _10195_/B _10195_/C vssd1 vssd1 vccd1 vccd1 _10196_/A sky130_fd_sc_hd__and3_1
XFILLER_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13954_ _13953_/X _13952_/Y _14612_/A vssd1 vssd1 vccd1 vccd1 _13954_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12905_ _12903_/Y _12899_/C _12901_/X _12902_/Y vssd1 vssd1 vccd1 vccd1 _12906_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13885_ _16086_/Q _14988_/A _13885_/C vssd1 vssd1 vccd1 vccd1 _13895_/A sky130_fd_sc_hd__and3_1
XFILLER_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15624_ _15194_/Q _15624_/D vssd1 vssd1 vccd1 vccd1 _15624_/Q sky130_fd_sc_hd__dfxtp_1
X_12836_ _12851_/A _12836_/B _12836_/C vssd1 vssd1 vccd1 vccd1 _12837_/A sky130_fd_sc_hd__and3_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _15655_/CLK _15555_/D vssd1 vssd1 vccd1 vccd1 _15555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _13041_/A vssd1 vssd1 vccd1 vccd1 _12767_/X sky130_fd_sc_hd__buf_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14517_/A _14506_/B _14510_/A vssd1 vssd1 vccd1 vccd1 _16207_/D sky130_fd_sc_hd__nor3_1
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11718_ _11796_/A _11718_/B _11722_/B vssd1 vssd1 vccd1 vccd1 _15725_/D sky130_fd_sc_hd__nor3_1
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15486_ _15224_/Q _15486_/D vssd1 vssd1 vccd1 vccd1 _15486_/Q sky130_fd_sc_hd__dfxtp_2
X_12698_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12740_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14437_ _14442_/A _14436_/Y _14431_/B _14432_/C vssd1 vssd1 vccd1 vccd1 _14439_/B
+ sky130_fd_sc_hd__o211a_1
X_11649_ _15716_/Q _11655_/C _11472_/X vssd1 vssd1 vccd1 vccd1 _11649_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14368_ _14368_/A vssd1 vssd1 vccd1 vccd1 _14368_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16107_ _16367_/CLK _16107_/D vssd1 vssd1 vccd1 vccd1 _16107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13319_ _15984_/Q _13420_/B _13319_/C vssd1 vssd1 vccd1 vccd1 _13324_/A sky130_fd_sc_hd__and3_1
X_14299_ _16167_/Q _14474_/B _14299_/C vssd1 vssd1 vccd1 vccd1 _14307_/A sky130_fd_sc_hd__and3_1
XFILLER_143_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16038_ _16050_/CLK _16038_/D vssd1 vssd1 vccd1 vccd1 _16038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08860_ _15283_/Q _08867_/C _08625_/X vssd1 vssd1 vccd1 vccd1 _08860_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07811_ _15737_/Q _08056_/B vssd1 vssd1 vccd1 vccd1 _08059_/B sky130_fd_sc_hd__xnor2_2
X_08791_ _08811_/C vssd1 vssd1 vccd1 vccd1 _08823_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07742_ _15936_/Q vssd1 vssd1 vccd1 vccd1 _13097_/C sky130_fd_sc_hd__clkinv_4
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07673_ _10965_/C vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09412_ _15367_/Q _09411_/C _09180_/X vssd1 vssd1 vccd1 vccd1 _09413_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09343_ _09339_/X _09340_/Y _09342_/Y _09337_/C vssd1 vssd1 vccd1 vccd1 _09345_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_21_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09274_ _09288_/A _09274_/B _09274_/C vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__and3_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08225_ _08225_/A _08105_/A vssd1 vssd1 vccd1 vccd1 _08231_/B sky130_fd_sc_hd__or2b_1
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08156_ _15270_/Q _08156_/B vssd1 vssd1 vccd1 vccd1 _08156_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08087_ _15539_/Q vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__clkinv_2
XFILLER_122_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08989_ _15301_/Q _09047_/B _08989_/C vssd1 vssd1 vccd1 vccd1 _08989_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10951_ _10946_/X _10949_/Y _10950_/Y _10944_/C vssd1 vssd1 vccd1 vccd1 _10953_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_29_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ _16035_/Q vssd1 vssd1 vccd1 vccd1 _13675_/C sky130_fd_sc_hd__inv_2
X_10882_ _15597_/Q _10999_/B _10882_/C vssd1 vssd1 vccd1 vccd1 _10882_/X sky130_fd_sc_hd__and3_1
X_12621_ _12621_/A _12621_/B _12621_/C vssd1 vssd1 vccd1 vccd1 _12622_/A sky130_fd_sc_hd__and3_1
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15340_ _15368_/CLK _15340_/D vssd1 vssd1 vccd1 vccd1 _15340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _15859_/Q _12667_/B _12554_/C vssd1 vssd1 vccd1 vccd1 _12552_/X sky130_fd_sc_hd__and3_1
XFILLER_129_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ _11518_/C vssd1 vssd1 vccd1 vccd1 _11528_/C sky130_fd_sc_hd__clkbuf_1
X_15271_ _16352_/CLK _15271_/D vssd1 vssd1 vccd1 vccd1 _15271_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12483_ _15847_/Q _12593_/B _12492_/C vssd1 vssd1 vccd1 vccd1 _12488_/A sky130_fd_sc_hd__and3_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_14222_ _16150_/Q _14228_/C _14177_/X vssd1 vssd1 vccd1 vccd1 _14224_/B sky130_fd_sc_hd__a21oi_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11434_ _11434_/A _11434_/B vssd1 vssd1 vccd1 vccd1 _11435_/B sky130_fd_sc_hd__nor2_1
X_14153_ _14326_/A vssd1 vssd1 vccd1 vccd1 _14153_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11365_ _11365_/A _11365_/B _11365_/C vssd1 vssd1 vccd1 vccd1 _11366_/A sky130_fd_sc_hd__and3_1
X_13104_ _13105_/B _13105_/C _13105_/A vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__a21o_1
X_10316_ _10316_/A vssd1 vssd1 vccd1 vccd1 _15507_/D sky130_fd_sc_hd__clkbuf_1
X_14084_ _14123_/A _14084_/B _14084_/C vssd1 vssd1 vccd1 vccd1 _14085_/A sky130_fd_sc_hd__and3_1
X_11296_ _15661_/Q _11525_/B _11298_/C vssd1 vssd1 vccd1 vccd1 _11296_/X sky130_fd_sc_hd__and3_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _15942_/Q _15944_/Q _15943_/Q _12981_/X vssd1 vssd1 vccd1 vccd1 _15935_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_112_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10247_ _15498_/Q _10363_/B _10247_/C vssd1 vssd1 vccd1 vccd1 _10247_/X sky130_fd_sc_hd__and3_1
XFILLER_79_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10178_ _10191_/C vssd1 vssd1 vccd1 vccd1 _10199_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14986_ _14986_/A vssd1 vssd1 vccd1 vccd1 _16316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13937_ _16093_/Q _14117_/B _13937_/C vssd1 vssd1 vccd1 vccd1 _13942_/A sky130_fd_sc_hd__and3_1
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13868_ _13868_/A vssd1 vssd1 vccd1 vccd1 _13980_/A sky130_fd_sc_hd__buf_2
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15607_ _15194_/Q _15607_/D vssd1 vssd1 vccd1 vccd1 _15607_/Q sky130_fd_sc_hd__dfxtp_1
X_12819_ _15899_/Q vssd1 vssd1 vccd1 vccd1 _12832_/C sky130_fd_sc_hd__inv_2
X_13799_ _16069_/Q _14093_/B _13799_/C vssd1 vssd1 vccd1 vccd1 _13808_/A sky130_fd_sc_hd__and3_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15538_ _15655_/CLK _15538_/D vssd1 vssd1 vccd1 vccd1 _15538_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15469_ _15483_/CLK _15469_/D vssd1 vssd1 vccd1 vccd1 _15469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08010_ _08010_/A _08010_/B vssd1 vssd1 vccd1 vccd1 _08011_/B sky130_fd_sc_hd__and2_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09961_ _09955_/B _09956_/C _09958_/X _09959_/Y vssd1 vssd1 vccd1 vccd1 _09962_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08912_ _15291_/Q _09146_/B _08919_/C vssd1 vssd1 vccd1 vccd1 _08916_/B sky130_fd_sc_hd__nand3_1
X_09892_ _09925_/C vssd1 vssd1 vccd1 vccd1 _09931_/C sky130_fd_sc_hd__clkbuf_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _15296_/Q _15295_/Q _15294_/Q _08604_/X vssd1 vssd1 vccd1 vccd1 _15279_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08774_ _08774_/A _08774_/B _08778_/B vssd1 vssd1 vccd1 vccd1 _15267_/D sky130_fd_sc_hd__nor3_1
XFILLER_84_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07725_ _15279_/Q _15261_/Q vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07656_ _13640_/A vssd1 vssd1 vccd1 vccd1 _14993_/A sky130_fd_sc_hd__buf_4
XFILLER_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09326_ _15355_/Q _09496_/B _09326_/C vssd1 vssd1 vccd1 vccd1 _09326_/X sky130_fd_sc_hd__and3_1
X_09257_ _09270_/C vssd1 vssd1 vccd1 vccd1 _09278_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08208_ _08014_/A _08014_/B _08206_/X _08207_/Y vssd1 vssd1 vccd1 vccd1 _08209_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09188_ input8/X vssd1 vssd1 vccd1 vccd1 _10341_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08139_ _08139_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__xnor2_4
XFILLER_146_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11150_ _11267_/A vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10101_ _15474_/Q _10106_/C _09981_/X vssd1 vssd1 vccd1 vccd1 _10101_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11081_ _12230_/A vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10032_ _15463_/Q _10150_/B _10037_/C vssd1 vssd1 vccd1 vccd1 _10032_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14840_ _14840_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14842_/A sky130_fd_sc_hd__or2_1
XFILLER_124_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14771_ _14771_/A _14771_/B vssd1 vssd1 vccd1 vccd1 _16267_/D sky130_fd_sc_hd__nor2_1
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11983_ _11983_/A vssd1 vssd1 vccd1 vccd1 _15767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13722_ _13666_/X _13718_/C _13721_/Y vssd1 vssd1 vccd1 vccd1 _16052_/D sky130_fd_sc_hd__a21oi_1
X_10934_ _15605_/Q _10939_/B _10933_/X vssd1 vssd1 vccd1 vccd1 _10936_/C sky130_fd_sc_hd__a21o_1
XFILLER_17_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ _13730_/A _13653_/B _13658_/B vssd1 vssd1 vccd1 vccd1 _16040_/D sky130_fd_sc_hd__nor3_1
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ _10902_/A _10865_/B _10865_/C vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__and3_1
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12604_ _12598_/B _12599_/C _12601_/X _12602_/Y vssd1 vssd1 vccd1 vccd1 _12605_/C
+ sky130_fd_sc_hd__a211o_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _16031_/Q _13583_/C _13534_/X vssd1 vssd1 vccd1 vccd1 _13584_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10796_ _10794_/Y _10789_/C _10801_/A _10793_/Y vssd1 vssd1 vccd1 vccd1 _10801_/B
+ sky130_fd_sc_hd__a211oi_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15323_ _15368_/CLK _15323_/D vssd1 vssd1 vccd1 vccd1 _15323_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _12554_/C vssd1 vssd1 vccd1 vccd1 _12568_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15254_ _15254_/CLK _15254_/D vssd1 vssd1 vccd1 vccd1 _15254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12466_ _12466_/A _12466_/B vssd1 vssd1 vccd1 vccd1 _12471_/C sky130_fd_sc_hd__nor2_1
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14205_ _14216_/C vssd1 vssd1 vccd1 vccd1 _14228_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11417_ _15679_/Q _11650_/B _11423_/C vssd1 vssd1 vccd1 vccd1 _11417_/Y sky130_fd_sc_hd__nand3_1
X_15185_ _15001_/A _15178_/A _15181_/B _15184_/Y vssd1 vssd1 vccd1 vccd1 _16364_/D
+ sky130_fd_sc_hd__o31a_1
X_12397_ _12397_/A vssd1 vssd1 vccd1 vccd1 _15832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14136_ _14133_/B _14132_/Y _14133_/A vssd1 vssd1 vccd1 vccd1 _14136_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_4_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ _15669_/Q _11355_/C _11230_/X vssd1 vssd1 vccd1 vccd1 _11348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14067_ _14080_/C vssd1 vssd1 vccd1 vccd1 _14093_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11279_ _15658_/Q _11317_/C _11047_/X vssd1 vssd1 vccd1 vccd1 _11281_/B sky130_fd_sc_hd__a21oi_1
XFILLER_140_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13018_ _15932_/Q _13018_/B _13022_/C vssd1 vssd1 vccd1 vccd1 _13018_/Y sky130_fd_sc_hd__nand3_1
XFILLER_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14969_ _14969_/A _14969_/B vssd1 vssd1 vccd1 vccd1 _16312_/D sky130_fd_sc_hd__nor2_1
XFILLER_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08490_ _08490_/A vssd1 vssd1 vccd1 vccd1 _15227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ _15321_/Q _09117_/C _08873_/X vssd1 vssd1 vccd1 vccd1 _09111_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09042_ _09036_/B _09037_/C _09039_/X _09040_/Y vssd1 vssd1 vccd1 vccd1 _09043_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_136_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09944_ _10388_/A vssd1 vssd1 vccd1 vccd1 _10064_/A sky130_fd_sc_hd__buf_2
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09875_ _15439_/Q _09874_/C _09755_/X vssd1 vssd1 vccd1 vccd1 _09876_/B sky130_fd_sc_hd__a21oi_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _15276_/Q _08947_/B _08831_/C vssd1 vssd1 vccd1 vccd1 _08826_/Y sky130_fd_sc_hd__nand3_1
XFILLER_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08757_ _08757_/A vssd1 vssd1 vccd1 vccd1 _15265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _12639_/A vssd1 vssd1 vccd1 vccd1 _12758_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08688_ _08686_/X _08687_/Y _08682_/B _08683_/C vssd1 vssd1 vccd1 vccd1 _08690_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_54_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _15017_/A _07639_/B _07639_/C vssd1 vssd1 vccd1 vccd1 _07640_/A sky130_fd_sc_hd__and3_1
XFILLER_26_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ _10651_/B _10651_/C _10651_/A vssd1 vssd1 vccd1 vccd1 _10652_/B sky130_fd_sc_hd__a21o_1
X_09309_ _09345_/A _09309_/B _09309_/C vssd1 vssd1 vccd1 vccd1 _09310_/A sky130_fd_sc_hd__and3_1
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10581_ _15556_/Q _15555_/Q _15554_/Q _10409_/X vssd1 vssd1 vccd1 vccd1 _15548_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12320_ _12314_/B _12315_/C _12317_/X _12318_/Y vssd1 vssd1 vccd1 vccd1 _12321_/C
+ sky130_fd_sc_hd__a211o_1
X_12251_ _12270_/C vssd1 vssd1 vccd1 vccd1 _12284_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ _11202_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11203_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _12182_/A _12182_/B vssd1 vssd1 vccd1 vccd1 _12187_/C sky130_fd_sc_hd__nor2_1
XFILLER_123_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11133_ _11133_/A _11133_/B _11133_/C vssd1 vssd1 vccd1 vccd1 _11134_/A sky130_fd_sc_hd__and3_1
XFILLER_123_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11064_ _15625_/Q _11236_/B _11066_/C vssd1 vssd1 vccd1 vccd1 _11064_/X sky130_fd_sc_hd__and3_1
X_15941_ _15196_/Q _15941_/D vssd1 vssd1 vccd1 vccd1 _15941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10015_ _10015_/A vssd1 vssd1 vccd1 vccd1 _15460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15872_ _15899_/CLK _15872_/D vssd1 vssd1 vccd1 vccd1 _15872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14823_ _15021_/A vssd1 vssd1 vccd1 vccd1 _14977_/B sky130_fd_sc_hd__buf_2
XFILLER_17_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11966_ _11978_/C vssd1 vssd1 vccd1 vccd1 _11986_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14754_ _14825_/A _14754_/B _14758_/B vssd1 vssd1 vccd1 vccd1 _16263_/D sky130_fd_sc_hd__nor3_1
XFILLER_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _10915_/A _10915_/B _10916_/X vssd1 vssd1 vccd1 vccd1 _15600_/D sky130_fd_sc_hd__a21oi_1
X_13705_ _13703_/Y _13698_/C _13711_/A _13702_/Y vssd1 vssd1 vccd1 vccd1 _13711_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_17_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14685_ _14883_/A vssd1 vssd1 vccd1 vccd1 _14847_/A sky130_fd_sc_hd__buf_2
X_11897_ _11895_/A _11895_/B _11896_/X vssd1 vssd1 vccd1 vccd1 _15753_/D sky130_fd_sc_hd__a21oi_1
XFILLER_149_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13636_ _13634_/X _13635_/Y _13631_/B _13632_/C vssd1 vssd1 vccd1 vccd1 _13638_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10848_ _11137_/A vssd1 vssd1 vccd1 vccd1 _10848_/X sky130_fd_sc_hd__buf_2
XFILLER_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16355_ _16358_/CLK _16355_/D vssd1 vssd1 vccd1 vccd1 _16355_/Q sky130_fd_sc_hd__dfxtp_1
X_13567_ _13412_/X _13564_/C _13566_/Y vssd1 vssd1 vccd1 vccd1 _16025_/D sky130_fd_sc_hd__a21oi_1
X_10779_ _10776_/X _10777_/Y _10778_/Y _10774_/C vssd1 vssd1 vccd1 vccd1 _10781_/B
+ sky130_fd_sc_hd__o211ai_1
X_15306_ _15339_/CLK _15306_/D vssd1 vssd1 vccd1 vccd1 _15306_/Q sky130_fd_sc_hd__dfxtp_4
X_12518_ _12518_/A _12518_/B _12522_/B vssd1 vssd1 vccd1 vccd1 _15851_/D sky130_fd_sc_hd__nor3_1
XFILLER_118_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16286_ _16321_/CLK _16286_/D vssd1 vssd1 vccd1 vccd1 _16286_/Q sky130_fd_sc_hd__dfxtp_1
X_13498_ _16015_/Q _13648_/B _13498_/C vssd1 vssd1 vccd1 vccd1 _13507_/A sky130_fd_sc_hd__and3_1
XFILLER_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15237_ _15926_/CLK _15237_/D vssd1 vssd1 vccd1 vccd1 _15237_/Q sky130_fd_sc_hd__dfxtp_1
X_12449_ _15842_/Q _12675_/B _12456_/C vssd1 vssd1 vccd1 vccd1 _12449_/X sky130_fd_sc_hd__and3_1
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15168_ _15168_/A _15168_/B _15168_/C vssd1 vssd1 vccd1 vccd1 _15169_/C sky130_fd_sc_hd__nand3_1
XFILLER_114_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14119_ _16130_/Q _14249_/B _14125_/C vssd1 vssd1 vccd1 vccd1 _14122_/B sky130_fd_sc_hd__nand3_1
X_15099_ _15099_/A _15099_/B _15099_/C vssd1 vssd1 vccd1 vccd1 _15100_/C sky130_fd_sc_hd__nand3_1
X_07990_ _13729_/C _07857_/B _07989_/X vssd1 vssd1 vccd1 vccd1 _08002_/A sky130_fd_sc_hd__o21ai_4
XFILLER_140_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09660_ _09680_/C vssd1 vssd1 vccd1 vccd1 _09692_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08611_ _08611_/A _08611_/B _08619_/A vssd1 vssd1 vccd1 vccd1 _15244_/D sky130_fd_sc_hd__nor3_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09591_ _09589_/A _09589_/B _09590_/X vssd1 vssd1 vccd1 vccd1 _15393_/D sky130_fd_sc_hd__a21oi_1
X_08542_ _08540_/B _08540_/C _08541_/X vssd1 vssd1 vccd1 vccd1 _08543_/C sky130_fd_sc_hd__o21ai_1
XFILLER_35_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08473_ _08944_/A vssd1 vssd1 vccd1 vccd1 _08611_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _09039_/C vssd1 vssd1 vccd1 vccd1 _09047_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _15446_/Q _10102_/B _09931_/C vssd1 vssd1 vccd1 vccd1 _09927_/Y sky130_fd_sc_hd__nand3_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09858_ _09865_/A _09858_/B _09858_/C vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__and3_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08809_ _15275_/Q _08811_/C _08634_/X vssd1 vssd1 vccd1 vccd1 _08809_/Y sky130_fd_sc_hd__a21oi_1
X_09789_ _09781_/B _09782_/C _09784_/X _09787_/Y vssd1 vssd1 vccd1 vccd1 _09790_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_46_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _15743_/Q _11827_/C _11760_/X vssd1 vssd1 vccd1 vccd1 _11820_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _15733_/Q _11811_/B _11754_/C vssd1 vssd1 vccd1 vccd1 _11751_/X sky130_fd_sc_hd__and3_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15395_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _10722_/C vssd1 vssd1 vccd1 vccd1 _10734_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _14471_/B _14471_/C _14471_/A vssd1 vssd1 vccd1 vccd1 _14472_/B sky130_fd_sc_hd__a21o_1
X_11682_ _11796_/A _11682_/B _11686_/A vssd1 vssd1 vccd1 vccd1 _15720_/D sky130_fd_sc_hd__nor3_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13421_ _13476_/A _13421_/B _13427_/A vssd1 vssd1 vccd1 vccd1 _16000_/D sky130_fd_sc_hd__nor3_1
X_10633_ _11783_/A vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__buf_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16140_ _16143_/CLK _16140_/D vssd1 vssd1 vccd1 vccd1 _16140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _13352_/A _13352_/B vssd1 vssd1 vccd1 vccd1 _13353_/B sky130_fd_sc_hd__nor2_1
X_10564_ _15545_/Q _10681_/B _10569_/C vssd1 vssd1 vccd1 vccd1 _10564_/Y sky130_fd_sc_hd__nand3_1
X_12303_ _15826_/Q _15825_/Q _15824_/Q _12134_/X vssd1 vssd1 vccd1 vccd1 _15818_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_6_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16071_ _16123_/CLK _16071_/D vssd1 vssd1 vccd1 vccd1 _16071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13283_ _13283_/A vssd1 vssd1 vccd1 vccd1 _13339_/A sky130_fd_sc_hd__clkbuf_2
X_10495_ _10503_/A _10495_/B _10495_/C vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__and3_1
X_15022_ _16328_/Q _15163_/B _15024_/C vssd1 vssd1 vccd1 vccd1 _15027_/A sky130_fd_sc_hd__and3_1
XFILLER_5_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12234_ _12234_/A _12234_/B _12238_/B vssd1 vssd1 vccd1 vccd1 _15806_/D sky130_fd_sc_hd__nor3_1
XFILLER_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12165_ _15797_/Q _12391_/B _12172_/C vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__and3_1
XFILLER_146_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ _11110_/B _11111_/C _11113_/X _11114_/Y vssd1 vssd1 vccd1 vccd1 _11117_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12096_ _12089_/B _12090_/C _12092_/X _12094_/Y vssd1 vssd1 vccd1 vccd1 _12097_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_110_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11047_ _11624_/A vssd1 vssd1 vccd1 vccd1 _11047_/X sky130_fd_sc_hd__buf_2
X_15924_ _07603_/A _15924_/D vssd1 vssd1 vccd1 vccd1 _15924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 reset vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_4
XFILLER_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15855_ _07603_/A _15855_/D vssd1 vssd1 vccd1 vccd1 _15855_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14806_ _14806_/A vssd1 vssd1 vccd1 vccd1 _14963_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15786_ _15794_/CLK _15786_/D vssd1 vssd1 vccd1 vccd1 _15786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12998_ _12996_/X _12997_/Y _12993_/B _12994_/C vssd1 vssd1 vccd1 vccd1 _13000_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_92_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14737_ _14936_/A vssd1 vssd1 vccd1 vccd1 _14825_/A sky130_fd_sc_hd__clkbuf_2
X_11949_ _11949_/A _11949_/B _11953_/B vssd1 vssd1 vccd1 vccd1 _15761_/D sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_71_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15301_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14668_ _14668_/A _14668_/B _14668_/C vssd1 vssd1 vccd1 vccd1 _14669_/C sky130_fd_sc_hd__nand3_1
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _13412_/X _13615_/C _13618_/Y vssd1 vssd1 vccd1 vccd1 _16034_/D sky130_fd_sc_hd__a21oi_1
X_14599_ _16231_/Q _14605_/C _13293_/B vssd1 vssd1 vccd1 vccd1 _14601_/B sky130_fd_sc_hd__a21oi_1
XFILLER_146_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16338_ _16359_/CLK _16338_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16269_ _16321_/CLK _16269_/D vssd1 vssd1 vccd1 vccd1 _16269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07973_ _07973_/A _07973_/B vssd1 vssd1 vccd1 vccd1 _07974_/B sky130_fd_sc_hd__and2_1
XFILLER_141_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ _15421_/Q _15420_/Q _15419_/Q _09541_/X vssd1 vssd1 vccd1 vccd1 _15413_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_68_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09643_ _09643_/A _09643_/B _09647_/B vssd1 vssd1 vccd1 vccd1 _15401_/D sky130_fd_sc_hd__nor3_1
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09574_ _09572_/Y _09568_/C _09570_/X _09571_/Y vssd1 vssd1 vccd1 vccd1 _09575_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08525_ _15232_/Q _08532_/C _08524_/X vssd1 vssd1 vccd1 vccd1 _08525_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16358_/CLK sky130_fd_sc_hd__clkbuf_16
X_08456_ _15017_/A _08456_/B _08456_/C vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__and3_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08387_ _08387_/A _08387_/B vssd1 vssd1 vccd1 vccd1 _08388_/B sky130_fd_sc_hd__nor2_2
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09008_ hold29/A _09067_/B _09008_/C vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__and3_1
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ _10280_/A _10280_/B vssd1 vssd1 vccd1 vccd1 _10284_/C sky130_fd_sc_hd__nor2_1
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13970_ _14413_/A _15013_/A _13964_/B _13969_/X vssd1 vssd1 vccd1 vccd1 _13971_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12959_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15640_ _15655_/CLK _15640_/D vssd1 vssd1 vccd1 vccd1 _15640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12852_ _12852_/A vssd1 vssd1 vccd1 vccd1 _15904_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11803_ _11803_/A vssd1 vssd1 vccd1 vccd1 _15739_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _15655_/CLK _15571_/D vssd1 vssd1 vccd1 vccd1 _15571_/Q sky130_fd_sc_hd__dfxtp_1
X_12783_ _12783_/A vssd1 vssd1 vccd1 vccd1 _15893_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16283_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _11754_/C vssd1 vssd1 vccd1 vccd1 _11767_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14522_ _14521_/X _14520_/Y _14648_/A vssd1 vssd1 vccd1 vccd1 _14522_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11665_/A _11665_/B vssd1 vssd1 vccd1 vccd1 _11666_/B sky130_fd_sc_hd__nor2_1
X_14453_ _14532_/A _14453_/B vssd1 vssd1 vccd1 vccd1 _14454_/B sky130_fd_sc_hd__and2_1
X_10616_ _10616_/A vssd1 vssd1 vccd1 vccd1 _15553_/D sky130_fd_sc_hd__clkbuf_1
X_13404_ _13404_/A _13404_/B vssd1 vssd1 vccd1 vccd1 _13405_/B sky130_fd_sc_hd__nor2_1
X_14384_ _16184_/Q _14389_/C _14250_/X vssd1 vssd1 vccd1 vccd1 _14386_/C sky130_fd_sc_hd__a21o_1
X_11596_ _11594_/Y _11588_/C _11592_/X _11593_/Y vssd1 vssd1 vccd1 vccd1 _11597_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16123_ _16123_/CLK _16123_/D vssd1 vssd1 vccd1 vccd1 _16123_/Q sky130_fd_sc_hd__dfxtp_1
X_13335_ _14593_/B vssd1 vssd1 vccd1 vccd1 _13543_/B sky130_fd_sc_hd__clkbuf_4
X_10547_ _15544_/Q _10549_/C _10373_/X vssd1 vssd1 vccd1 vccd1 _10547_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16054_ _16075_/CLK _16054_/D vssd1 vssd1 vccd1 vccd1 _16054_/Q sky130_fd_sc_hd__dfxtp_2
X_13266_ _15975_/Q _13420_/B _13266_/C vssd1 vssd1 vccd1 vccd1 _13272_/A sky130_fd_sc_hd__and3_1
X_10478_ _15533_/Q _10590_/B _10484_/C vssd1 vssd1 vccd1 vccd1 _10481_/B sky130_fd_sc_hd__nand3_1
X_12217_ _12214_/X _12215_/Y _12216_/Y _12212_/C vssd1 vssd1 vccd1 vccd1 _12219_/B
+ sky130_fd_sc_hd__o211ai_1
X_15005_ _15005_/A vssd1 vssd1 vccd1 vccd1 _15152_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13197_ _13197_/A _13197_/B vssd1 vssd1 vccd1 vccd1 _13198_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12148_ _12170_/A _12148_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12149_/A sky130_fd_sc_hd__and3_1
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12079_ _12102_/C vssd1 vssd1 vccd1 vccd1 _12115_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15907_ _15907_/CLK _15907_/D vssd1 vssd1 vccd1 vccd1 _15907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15838_ _07603_/A _15838_/D vssd1 vssd1 vccd1 vccd1 _15838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15769_ _15794_/CLK _15769_/D vssd1 vssd1 vccd1 vccd1 _15769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16204_/CLK sky130_fd_sc_hd__clkbuf_16
X_08310_ _08384_/A _08384_/C vssd1 vssd1 vccd1 vccd1 _08311_/B sky130_fd_sc_hd__xor2_1
X_09290_ _15349_/Q _09290_/B _09290_/C vssd1 vssd1 vccd1 vccd1 _09300_/A sky130_fd_sc_hd__and3_1
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08241_ _08241_/A _08241_/B vssd1 vssd1 vccd1 vccd1 _08249_/B sky130_fd_sc_hd__nand2_1
XANTENNA_14 _10751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _14541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_36 _13720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ _08163_/A _08163_/B _08171_/Y vssd1 vssd1 vccd1 vccd1 _08272_/A sky130_fd_sc_hd__a21bo_2
XFILLER_134_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07956_ _07887_/A _07887_/B _07886_/A vssd1 vssd1 vccd1 vccd1 _08195_/B sky130_fd_sc_hd__o21ai_2
X_07887_ _07887_/A _07887_/B vssd1 vssd1 vccd1 vccd1 _07888_/B sky130_fd_sc_hd__xor2_2
XFILLER_110_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09626_ _09635_/A _09626_/B _09626_/C vssd1 vssd1 vccd1 vccd1 _09627_/A sky130_fd_sc_hd__and3_1
XFILLER_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09557_ _15390_/Q _09784_/B _09557_/C vssd1 vssd1 vccd1 vccd1 _09557_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_35_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16367_/CLK sky130_fd_sc_hd__clkbuf_16
X_08508_ _08519_/A _08508_/B _08508_/C vssd1 vssd1 vccd1 vccd1 _08509_/A sky130_fd_sc_hd__and3_1
XFILLER_102_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09488_ _10065_/A vssd1 vssd1 vccd1 vccd1 _09721_/B sky130_fd_sc_hd__buf_2
XFILLER_24_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08439_ _08435_/Y _08437_/X _08438_/Y vssd1 vssd1 vccd1 vccd1 _15218_/D sky130_fd_sc_hd__a21oi_1
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11450_ _11509_/A _11450_/B _11454_/A vssd1 vssd1 vccd1 vccd1 _15684_/D sky130_fd_sc_hd__nor3_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ _10401_/A _10401_/B vssd1 vssd1 vccd1 vccd1 _10405_/C sky130_fd_sc_hd__nor2_1
X_11381_ _11555_/A vssd1 vssd1 vccd1 vccd1 _11420_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13120_ _14080_/B vssd1 vssd1 vccd1 vccd1 _14593_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ _10969_/A vssd1 vssd1 vccd1 vccd1 _11488_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_137_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13051_ _15940_/Q _13051_/B _13051_/C vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__and3_1
X_10263_ _15499_/Q _10441_/B _10268_/C vssd1 vssd1 vccd1 vccd1 _10263_/Y sky130_fd_sc_hd__nand3_1
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12002_ _15771_/Q _12007_/C _12001_/X vssd1 vssd1 vccd1 vccd1 _12002_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10194_ _10188_/B _10189_/C _10191_/X _10192_/Y vssd1 vssd1 vccd1 vccd1 _10195_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13953_ _13953_/A _13953_/B vssd1 vssd1 vccd1 vccd1 _13953_/X sky130_fd_sc_hd__or2_1
XFILLER_143_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _12901_/X _12902_/Y _12903_/Y _12899_/C vssd1 vssd1 vccd1 vccd1 _12906_/B
+ sky130_fd_sc_hd__o211ai_1
X_13884_ _14298_/A vssd1 vssd1 vccd1 vccd1 _14988_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15623_ _15194_/Q _15623_/D vssd1 vssd1 vccd1 vccd1 _15623_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _12829_/B _12830_/C _12832_/X _12833_/Y vssd1 vssd1 vccd1 vccd1 _12836_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _16119_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15655_/CLK _15554_/D vssd1 vssd1 vccd1 vccd1 _15554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12798_/C vssd1 vssd1 vccd1 vccd1 _12805_/C sky130_fd_sc_hd__clkbuf_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14505_ _16210_/Q _14546_/B _14505_/C vssd1 vssd1 vccd1 vccd1 _14510_/A sky130_fd_sc_hd__and3_1
X_11717_ _11715_/Y _11708_/C _11722_/A _11714_/Y vssd1 vssd1 vccd1 vccd1 _11722_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15485_ _15485_/CLK _15485_/D vssd1 vssd1 vccd1 vccd1 _15485_/Q sky130_fd_sc_hd__dfxtp_1
X_12697_ _12695_/A _12695_/B _12696_/X vssd1 vssd1 vccd1 vccd1 _15879_/D sky130_fd_sc_hd__a21oi_1
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11648_ _15716_/Q _11819_/B _11655_/C vssd1 vssd1 vccd1 vccd1 _11648_/X sky130_fd_sc_hd__and3_1
X_14436_ _16194_/Q _14435_/C _14300_/X vssd1 vssd1 vccd1 vccd1 _14436_/Y sky130_fd_sc_hd__a21oi_1
X_11579_ _11573_/B _11574_/C _11576_/X _11577_/Y vssd1 vssd1 vccd1 vccd1 _11580_/C
+ sky130_fd_sc_hd__a211o_1
X_14367_ _14190_/X _14365_/B _14366_/Y vssd1 vssd1 vccd1 vccd1 _16176_/D sky130_fd_sc_hd__o21a_1
X_16106_ _16222_/CLK _16106_/D vssd1 vssd1 vccd1 vccd1 _16106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13318_ _15984_/Q _13349_/C _13317_/X vssd1 vssd1 vccd1 vccd1 _13320_/B sky130_fd_sc_hd__a21oi_1
XFILLER_128_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14298_ _14298_/A vssd1 vssd1 vccd1 vccd1 _14474_/B sky130_fd_sc_hd__buf_2
XFILLER_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16037_ _16040_/CLK _16037_/D vssd1 vssd1 vccd1 vccd1 _16037_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13249_ _13249_/A _13249_/B vssd1 vssd1 vccd1 vccd1 _13252_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07810_ _15701_/Q _15719_/Q vssd1 vssd1 vccd1 vccd1 _08056_/B sky130_fd_sc_hd__xor2_2
XFILLER_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08790_ _08802_/C vssd1 vssd1 vccd1 vccd1 _08811_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_07741_ _15728_/Q _08136_/B vssd1 vssd1 vccd1 vccd1 _07757_/A sky130_fd_sc_hd__xnor2_4
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07672_ _07672_/A vssd1 vssd1 vccd1 vccd1 _10965_/C sky130_fd_sc_hd__buf_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09411_ _15367_/Q _09644_/B _09411_/C vssd1 vssd1 vccd1 vccd1 _09419_/B sky130_fd_sc_hd__and3_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _16050_/CLK sky130_fd_sc_hd__clkbuf_16
X_09342_ _15356_/Q _09572_/B _09348_/C vssd1 vssd1 vccd1 vccd1 _09342_/Y sky130_fd_sc_hd__nand3_1
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09273_ _09266_/B _09267_/C _09270_/X _09271_/Y vssd1 vssd1 vccd1 vccd1 _09274_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08224_ _08224_/A _08104_/A vssd1 vssd1 vccd1 vccd1 _08231_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08173_/A sky130_fd_sc_hd__xnor2_4
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08086_ _15557_/Q vssd1 vssd1 vccd1 vccd1 _10639_/A sky130_fd_sc_hd__inv_2
XFILLER_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08988_ _15302_/Q _08989_/C _08929_/X vssd1 vssd1 vccd1 vccd1 _08988_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07939_ _10700_/A _07939_/B vssd1 vssd1 vccd1 vccd1 _07942_/B sky130_fd_sc_hd__xnor2_1
XFILLER_91_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10950_ _15606_/Q _10950_/B _10950_/C vssd1 vssd1 vccd1 vccd1 _10950_/Y sky130_fd_sc_hd__nand3_1
XFILLER_113_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09609_ _15398_/Q _09721_/B _09615_/C vssd1 vssd1 vccd1 vccd1 _09612_/B sky130_fd_sc_hd__nand3_1
X_10881_ _10881_/A vssd1 vssd1 vccd1 vccd1 _15595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12620_ _12618_/Y _12613_/C _12615_/X _12617_/Y vssd1 vssd1 vccd1 vccd1 _12621_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _12551_/A vssd1 vssd1 vccd1 vccd1 _15857_/D sky130_fd_sc_hd__clkbuf_1
X_11502_ _11502_/A vssd1 vssd1 vccd1 vccd1 _11518_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15270_ _15282_/CLK _15270_/D vssd1 vssd1 vccd1 vccd1 _15270_/Q sky130_fd_sc_hd__dfxtp_1
X_12482_ _15847_/Q _12519_/C _12481_/X vssd1 vssd1 vccd1 vccd1 _12484_/B sky130_fd_sc_hd__a21oi_1
X_11433_ _11439_/B _11433_/B vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__or2_1
X_14221_ _16150_/Q _14221_/B _14228_/C vssd1 vssd1 vccd1 vccd1 _14224_/A sky130_fd_sc_hd__and3_1
XFILLER_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14152_ _14058_/X _14146_/B _14059_/X vssd1 vssd1 vccd1 vccd1 _14155_/A sky130_fd_sc_hd__a21oi_1
X_11364_ _11362_/Y _11358_/C _11360_/X _11361_/Y vssd1 vssd1 vccd1 vccd1 _11365_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10315_ _10323_/A _10315_/B _10315_/C vssd1 vssd1 vccd1 vccd1 _10316_/A sky130_fd_sc_hd__and3_1
X_13103_ _15949_/Q _13109_/C _14250_/A vssd1 vssd1 vccd1 vccd1 _13105_/C sky130_fd_sc_hd__a21o_1
X_14083_ _14077_/B _14078_/C _14080_/X _14081_/Y vssd1 vssd1 vccd1 vccd1 _14084_/C
+ sky130_fd_sc_hd__a211o_1
X_11295_ _11582_/A vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _13034_/A vssd1 vssd1 vccd1 vccd1 _15934_/D sky130_fd_sc_hd__clkbuf_1
X_10246_ _10246_/A vssd1 vssd1 vccd1 vccd1 _15496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10177_ _10177_/A vssd1 vssd1 vccd1 vccd1 _10191_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14985_ _15135_/A _14985_/B _14985_/C vssd1 vssd1 vccd1 vccd1 _14986_/A sky130_fd_sc_hd__and3_1
XFILLER_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13936_ _16093_/Q _13957_/C _13822_/X vssd1 vssd1 vccd1 vccd1 _13938_/B sky130_fd_sc_hd__a21oi_1
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13867_ _16097_/Q _16096_/Q _16095_/Q _13723_/X vssd1 vssd1 vccd1 vccd1 _16080_/D
+ sky130_fd_sc_hd__o31a_1
X_15606_ _15194_/Q _15606_/D vssd1 vssd1 vccd1 vccd1 _15606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12818_ _13239_/A vssd1 vssd1 vccd1 vccd1 _12934_/A sky130_fd_sc_hd__buf_2
X_13798_ _13798_/A vssd1 vssd1 vccd1 vccd1 _16066_/D sky130_fd_sc_hd__clkbuf_1
X_15537_ _15655_/CLK _15537_/D vssd1 vssd1 vccd1 vccd1 _15537_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _15889_/Q _12748_/C _12631_/X vssd1 vssd1 vccd1 vccd1 _12750_/B sky130_fd_sc_hd__a21oi_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15468_ _15483_/CLK _15468_/D vssd1 vssd1 vccd1 vccd1 _15468_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14419_ _14328_/X _14372_/X _14411_/B _14240_/X vssd1 vssd1 vccd1 vccd1 _14420_/B
+ sky130_fd_sc_hd__a31o_1
X_15399_ _15483_/CLK _15399_/D vssd1 vssd1 vccd1 vccd1 _15399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09960_ _09958_/X _09959_/Y _09955_/B _09956_/C vssd1 vssd1 vccd1 vccd1 _09962_/B
+ sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_6_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _15971_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08911_ _10065_/A vssd1 vssd1 vccd1 vccd1 _09146_/B sky130_fd_sc_hd__clkbuf_2
X_09891_ _09911_/C vssd1 vssd1 vccd1 vccd1 _09925_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08842_/A vssd1 vssd1 vccd1 vccd1 _15278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08771_/Y _08765_/C _08778_/A _08770_/Y vssd1 vssd1 vccd1 vccd1 _08778_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_84_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07724_ _15297_/Q vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__clkinv_2
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07655_ _12726_/A vssd1 vssd1 vccd1 vccd1 _13640_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09325_ _09325_/A vssd1 vssd1 vccd1 vccd1 _15353_/D sky130_fd_sc_hd__clkbuf_1
X_09256_ _09256_/A vssd1 vssd1 vccd1 vccd1 _09270_/C sky130_fd_sc_hd__clkbuf_2
X_08207_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08207_/Y sky130_fd_sc_hd__nor2_1
X_09187_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09233_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08138_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08139_/B sky130_fd_sc_hd__xor2_4
XFILLER_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08069_ _08069_/A _08069_/B vssd1 vssd1 vccd1 vccd1 _08226_/A sky130_fd_sc_hd__nand2_1
X_10100_ _15474_/Q _10155_/B _10100_/C vssd1 vssd1 vccd1 vccd1 _10109_/A sky130_fd_sc_hd__and3_1
X_11080_ _11080_/A vssd1 vssd1 vccd1 vccd1 _12230_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10031_ _15464_/Q _10037_/C _10030_/X vssd1 vssd1 vccd1 vccd1 _10031_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ _14694_/X _14768_/A _14695_/X vssd1 vssd1 vccd1 vccd1 _14771_/B sky130_fd_sc_hd__o21ai_1
X_11982_ _11997_/A _11982_/B _11982_/C vssd1 vssd1 vccd1 vccd1 _11983_/A sky130_fd_sc_hd__and3_1
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13721_ _13617_/X _13718_/C _13720_/X vssd1 vssd1 vccd1 vccd1 _13721_/Y sky130_fd_sc_hd__o21ai_1
X_10933_ _11222_/A vssd1 vssd1 vccd1 vccd1 _10933_/X sky130_fd_sc_hd__buf_2
XFILLER_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10864_ _10863_/B _10863_/C _10751_/X vssd1 vssd1 vccd1 vccd1 _10865_/C sky130_fd_sc_hd__o21ai_1
X_13652_ _13650_/Y _13646_/C _13658_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13658_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12603_ _12601_/X _12602_/Y _12598_/B _12599_/C vssd1 vssd1 vccd1 vccd1 _12605_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _16031_/Q _13738_/B _13583_/C vssd1 vssd1 vccd1 vccd1 _13583_/X sky130_fd_sc_hd__and3_1
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10795_ _10801_/A _10793_/Y _10794_/Y _10789_/C vssd1 vssd1 vccd1 vccd1 _10797_/B
+ sky130_fd_sc_hd__o211a_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _15322_/CLK _15322_/D vssd1 vssd1 vccd1 vccd1 _15322_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12546_/C vssd1 vssd1 vccd1 vccd1 _12554_/C sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15253_ _15254_/CLK _15253_/D vssd1 vssd1 vccd1 vccd1 _15253_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12465_ _12465_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12466_/B sky130_fd_sc_hd__nor2_1
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14204_ _14207_/C vssd1 vssd1 vccd1 vccd1 _14216_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_144_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11416_ _12277_/A vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__buf_2
X_12396_ _12396_/A _12396_/B _12396_/C vssd1 vssd1 vccd1 vccd1 _12397_/A sky130_fd_sc_hd__and3_1
X_15184_ _15184_/A _15189_/C vssd1 vssd1 vccd1 vccd1 _15184_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11347_ _15669_/Q _11576_/B _11347_/C vssd1 vssd1 vccd1 vccd1 _11347_/X sky130_fd_sc_hd__and3_1
X_14135_ _14133_/A _14133_/B _14132_/Y _14134_/Y vssd1 vssd1 vccd1 vccd1 _16129_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_113_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ _11311_/C vssd1 vssd1 vccd1 vccd1 _11317_/C sky130_fd_sc_hd__clkbuf_2
X_14066_ _14071_/C vssd1 vssd1 vccd1 vccd1 _14080_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10229_ _10228_/B _10228_/C _10172_/X vssd1 vssd1 vccd1 vccd1 _10230_/C sky130_fd_sc_hd__o21ai_1
X_13017_ _15933_/Q _13022_/C _12855_/X vssd1 vssd1 vccd1 vccd1 _13017_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14968_ _14892_/X _14966_/A _14893_/X vssd1 vssd1 vccd1 vccd1 _14969_/B sky130_fd_sc_hd__o21ai_1
X_13919_ _13919_/A vssd1 vssd1 vccd1 vccd1 _13920_/A sky130_fd_sc_hd__buf_2
XFILLER_35_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14899_ hold28/X vssd1 vssd1 vccd1 vccd1 _14905_/C sky130_fd_sc_hd__inv_2
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ _15321_/Q _09165_/B _09117_/C vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__and3_1
XFILLER_148_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09041_ _09039_/X _09040_/Y _09036_/B _09037_/C vssd1 vssd1 vccd1 vccd1 _09043_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ _15457_/Q _15456_/Q _15455_/Q _09831_/X vssd1 vssd1 vccd1 vccd1 _15449_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09874_ _15439_/Q _09931_/B _09874_/C vssd1 vssd1 vccd1 vccd1 _09883_/B sky130_fd_sc_hd__and3_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08825_ _15277_/Q _08831_/C _08824_/X vssd1 vssd1 vccd1 vccd1 _08825_/Y sky130_fd_sc_hd__a21oi_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08756_ _08765_/A _08756_/B _08756_/C vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__and3_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07707_ _14814_/A vssd1 vssd1 vccd1 vccd1 _07707_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _15256_/Q _08694_/C _08625_/X vssd1 vssd1 vccd1 vccd1 _08687_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _07638_/A _07638_/B _07638_/C vssd1 vssd1 vccd1 vccd1 _07639_/C sky130_fd_sc_hd__nand3_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09308_ _09306_/B _09306_/C _09307_/X vssd1 vssd1 vccd1 vccd1 _09309_/C sky130_fd_sc_hd__o21ai_1
X_10580_ _10580_/A vssd1 vssd1 vccd1 vccd1 _15547_/D sky130_fd_sc_hd__clkbuf_1
X_09239_ _09245_/A _09237_/Y _09238_/Y _09233_/C vssd1 vssd1 vccd1 vccd1 _09241_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _12262_/C vssd1 vssd1 vccd1 vccd1 _12270_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ _11208_/B _11201_/B vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__or2_1
XFILLER_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12181_ _12181_/A _12181_/B vssd1 vssd1 vccd1 vccd1 _12182_/B sky130_fd_sc_hd__nor2_1
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11132_ _11130_/Y _11124_/C _11126_/X _11127_/Y vssd1 vssd1 vccd1 vccd1 _11133_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11063_ _11063_/A vssd1 vssd1 vccd1 vccd1 _15623_/D sky130_fd_sc_hd__clkbuf_1
X_15940_ _15196_/Q _15940_/D vssd1 vssd1 vccd1 vccd1 _15940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10014_ _10035_/A _10014_/B _10014_/C vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__and3_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15871_ _15907_/CLK _15871_/D vssd1 vssd1 vccd1 vccd1 _15871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14822_ _16283_/Q _14838_/C _14702_/X vssd1 vssd1 vccd1 vccd1 _14825_/B sky130_fd_sc_hd__a21oi_1
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14753_ _14747_/B _14748_/C _14758_/A _14751_/Y vssd1 vssd1 vccd1 vccd1 _14758_/B
+ sky130_fd_sc_hd__a211oi_1
X_11965_ _15764_/Q vssd1 vssd1 vccd1 vccd1 _11978_/C sky130_fd_sc_hd__inv_2
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13704_ _13711_/A _13702_/Y _13703_/Y _13698_/C vssd1 vssd1 vccd1 vccd1 _13706_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _10916_/A _10920_/C vssd1 vssd1 vccd1 vccd1 _10916_/X sky130_fd_sc_hd__or2_1
X_14684_ _14682_/A _14682_/B _14683_/X vssd1 vssd1 vccd1 vccd1 _16246_/D sky130_fd_sc_hd__a21oi_1
X_11896_ _12068_/A _11901_/C vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__or2_1
X_13635_ _16040_/Q _13634_/C _13534_/X vssd1 vssd1 vccd1 vccd1 _13635_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10847_ _15591_/Q _11078_/B _10847_/C vssd1 vssd1 vccd1 vccd1 _10858_/A sky130_fd_sc_hd__and3_1
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16354_ _16358_/CLK _16354_/D vssd1 vssd1 vccd1 vccd1 _16354_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13566_ _13362_/X _13564_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13566_/Y sky130_fd_sc_hd__o21ai_1
X_10778_ _15579_/Q _10778_/B _10778_/C vssd1 vssd1 vccd1 vccd1 _10778_/Y sky130_fd_sc_hd__nand3_1
XFILLER_9_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15305_ _15359_/CLK _15305_/D vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
X_12517_ _12515_/Y _12510_/C _12522_/A _12513_/Y vssd1 vssd1 vccd1 vccd1 _12522_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16285_ _16321_/CLK _16285_/D vssd1 vssd1 vccd1 vccd1 _16285_/Q sky130_fd_sc_hd__dfxtp_1
X_13497_ _13868_/A vssd1 vssd1 vccd1 vccd1 _13604_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15236_ _15351_/CLK _15236_/D vssd1 vssd1 vccd1 vccd1 _15236_/Q sky130_fd_sc_hd__dfxtp_1
X_12448_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__buf_2
XFILLER_126_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15167_ _15168_/B _15168_/C _15168_/A vssd1 vssd1 vccd1 vccd1 _15169_/B sky130_fd_sc_hd__a21o_1
XFILLER_126_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ _12376_/X _12378_/Y _12373_/B _12374_/C vssd1 vssd1 vccd1 vccd1 _12381_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_141_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14118_ _14208_/A _14118_/B _14122_/A vssd1 vssd1 vccd1 vccd1 _16126_/D sky130_fd_sc_hd__nor3_1
XFILLER_140_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15098_ _15099_/B _15099_/C _15099_/A vssd1 vssd1 vccd1 vccd1 _15100_/B sky130_fd_sc_hd__a21o_1
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14049_ _14316_/A vssd1 vssd1 vccd1 vccd1 _14049_/X sky130_fd_sc_hd__buf_2
XFILLER_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ _15245_/Q _08794_/B _08610_/C vssd1 vssd1 vccd1 vccd1 _08619_/A sky130_fd_sc_hd__and3_1
X_09590_ _09760_/A _09594_/C vssd1 vssd1 vccd1 vccd1 _09590_/X sky130_fd_sc_hd__or2_1
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08541_ _12758_/A vssd1 vssd1 vccd1 vccd1 _08541_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08472_ _15242_/Q _15241_/Q _15240_/Q _07608_/X vssd1 vssd1 vccd1 vccd1 _15225_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09024_ _09024_/A vssd1 vssd1 vccd1 vccd1 _09039_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09926_ _15447_/Q _09931_/C _09693_/X vssd1 vssd1 vccd1 vccd1 _09926_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09857_ _09855_/Y _09851_/C _09853_/X _09854_/Y vssd1 vssd1 vccd1 vccd1 _09858_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08808_ _15275_/Q _08865_/B _08811_/C vssd1 vssd1 vccd1 vccd1 _08808_/X sky130_fd_sc_hd__and3_1
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09788_ _09784_/X _09787_/Y _09781_/B _09782_/C vssd1 vssd1 vccd1 vccd1 _09790_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _15264_/Q _08853_/B _08745_/C vssd1 vssd1 vccd1 vccd1 _08742_/B sky130_fd_sc_hd__nand3_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11750_/A vssd1 vssd1 vccd1 vccd1 _15731_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _10714_/C vssd1 vssd1 vccd1 vccd1 _10722_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _15721_/Q _11737_/B _11689_/C vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__and3_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13420_ _16002_/Q _13420_/B _13420_/C vssd1 vssd1 vccd1 vccd1 _13427_/A sky130_fd_sc_hd__and3_1
X_10632_ input8/X vssd1 vssd1 vccd1 vccd1 _11783_/A sky130_fd_sc_hd__buf_2
X_10563_ _15546_/Q _10569_/C _10562_/X vssd1 vssd1 vccd1 vccd1 _10563_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13351_ _13358_/B _13351_/B vssd1 vssd1 vccd1 vccd1 _13353_/A sky130_fd_sc_hd__or2_1
XFILLER_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ _12302_/A vssd1 vssd1 vccd1 vccd1 _15817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16070_ _16124_/CLK _16070_/D vssd1 vssd1 vccd1 vccd1 _16070_/Q sky130_fd_sc_hd__dfxtp_1
X_10494_ _10492_/Y _10488_/C _10490_/X _10491_/Y vssd1 vssd1 vccd1 vccd1 _10495_/C
+ sky130_fd_sc_hd__a211o_1
X_13282_ _13282_/A vssd1 vssd1 vccd1 vccd1 _15975_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15021_ _15021_/A vssd1 vssd1 vccd1 vccd1 _15163_/B sky130_fd_sc_hd__buf_2
X_12233_ _12231_/Y _12226_/C _12238_/A _12229_/Y vssd1 vssd1 vccd1 vccd1 _12238_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_107_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12164_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12391_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_111_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11115_ _11113_/X _11114_/Y _11110_/B _11111_/C vssd1 vssd1 vccd1 vccd1 _11117_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12095_ _12092_/X _12094_/Y _12089_/B _12090_/C vssd1 vssd1 vccd1 vccd1 _12097_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11046_ _11078_/C vssd1 vssd1 vccd1 vccd1 _11086_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15923_ _15196_/Q _15923_/D vssd1 vssd1 vccd1 vccd1 _15923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15854_ _15971_/CLK _15854_/D vssd1 vssd1 vccd1 vccd1 _15854_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14805_ _14802_/X _14797_/A _14800_/B _14804_/Y vssd1 vssd1 vccd1 vccd1 _16274_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15785_ _15794_/CLK _15785_/D vssd1 vssd1 vccd1 vccd1 _15785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12997_ _15930_/Q _13004_/C _13275_/A vssd1 vssd1 vccd1 vccd1 _12997_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14736_ hold13/X hold14/X hold12/X _14620_/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__o31a_1
X_11948_ _11946_/Y _11941_/C _11953_/A _11944_/Y vssd1 vssd1 vccd1 vccd1 _11953_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14667_ _14668_/B _14668_/C _14668_/A vssd1 vssd1 vccd1 vccd1 _14669_/B sky130_fd_sc_hd__a21o_1
X_11879_ _15752_/Q _11885_/C _11760_/X vssd1 vssd1 vccd1 vccd1 _11879_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13618_ _13617_/X _13615_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13618_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ _16231_/Q _14598_/B _14605_/C vssd1 vssd1 vccd1 vccd1 _14601_/A sky130_fd_sc_hd__and3_1
X_16337_ _16337_/CLK _16337_/D vssd1 vssd1 vccd1 vccd1 _16337_/Q sky130_fd_sc_hd__dfxtp_1
X_13549_ _16024_/Q _13554_/C _13342_/X vssd1 vssd1 vccd1 vccd1 _13549_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16268_ _16268_/CLK _16268_/D vssd1 vssd1 vccd1 vccd1 _16268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15219_ _16242_/CLK _15219_/D vssd1 vssd1 vccd1 vccd1 state1[4] sky130_fd_sc_hd__dfxtp_2
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16199_ _16247_/CLK _16199_/D vssd1 vssd1 vccd1 vccd1 _16199_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07972_ _07973_/A _07973_/B vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09711_ _09711_/A vssd1 vssd1 vccd1 vccd1 _15412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09642_ _09640_/Y _09635_/C _09647_/A _09639_/Y vssd1 vssd1 vccd1 vccd1 _09647_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_67_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09573_ _09570_/X _09571_/Y _09572_/Y _09568_/C vssd1 vssd1 vccd1 vccd1 _09575_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _09693_/A vssd1 vssd1 vccd1 vccd1 _08524_/X sky130_fd_sc_hd__buf_2
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08455_ _08465_/A _08453_/Y _08443_/A _08448_/A vssd1 vssd1 vccd1 vccd1 _08456_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08386_ _08386_/A _08386_/B _08386_/C vssd1 vssd1 vccd1 vccd1 _08387_/B sky130_fd_sc_hd__and3_1
XFILLER_149_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09007_ _09066_/A _09007_/B _09011_/B vssd1 vssd1 vccd1 vccd1 _15303_/D sky130_fd_sc_hd__nor3_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09909_ _15445_/Q _10022_/B _09911_/C vssd1 vssd1 vccd1 vccd1 _09909_/X sky130_fd_sc_hd__and3_1
XFILLER_76_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12920_ _12918_/A _12918_/B _12919_/X vssd1 vssd1 vccd1 vccd1 _15915_/D sky130_fd_sc_hd__a21oi_1
XFILLER_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _12851_/A _12851_/B _12851_/C vssd1 vssd1 vccd1 vccd1 _12852_/A sky130_fd_sc_hd__and3_1
XFILLER_92_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11802_ _11824_/A _11802_/B _11802_/C vssd1 vssd1 vccd1 vccd1 _11803_/A sky130_fd_sc_hd__and3_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15655_/CLK _15570_/D vssd1 vssd1 vccd1 vccd1 _15570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12796_/A _12782_/B _12782_/C vssd1 vssd1 vccd1 vccd1 _12783_/A sky130_fd_sc_hd__and3_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14521_/A _14521_/B vssd1 vssd1 vccd1 vccd1 _14521_/X sky130_fd_sc_hd__or2_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _11745_/C vssd1 vssd1 vccd1 vccd1 _11754_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14446_/Y _14447_/X _14449_/B vssd1 vssd1 vccd1 vccd1 _14453_/B sky130_fd_sc_hd__o21a_1
X_11664_ _11670_/B _11664_/B vssd1 vssd1 vccd1 vccd1 _11666_/A sky130_fd_sc_hd__or2_1
XFILLER_30_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ _13408_/B _13403_/B vssd1 vssd1 vccd1 vccd1 _13405_/A sky130_fd_sc_hd__or2_1
X_10615_ _10615_/A _10615_/B _10615_/C vssd1 vssd1 vccd1 vccd1 _10616_/A sky130_fd_sc_hd__and3_1
X_14383_ _16184_/Q _14468_/B _14389_/C vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__nand3_1
X_11595_ _11592_/X _11593_/Y _11594_/Y _11588_/C vssd1 vssd1 vccd1 vccd1 _11597_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16122_ _16123_/CLK _16122_/D vssd1 vssd1 vccd1 vccd1 _16122_/Q sky130_fd_sc_hd__dfxtp_1
X_13334_ _15987_/Q _13341_/C _13179_/X vssd1 vssd1 vccd1 vccd1 _13334_/Y sky130_fd_sc_hd__a21oi_1
X_10546_ _15544_/Q _10602_/B _10549_/C vssd1 vssd1 vccd1 vccd1 _10546_/X sky130_fd_sc_hd__and3_1
XFILLER_127_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16053_ _16075_/CLK _16053_/D vssd1 vssd1 vccd1 vccd1 _16053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13265_ _15975_/Q _13297_/C _13041_/X vssd1 vssd1 vccd1 vccd1 _13267_/B sky130_fd_sc_hd__a21oi_1
X_10477_ _10511_/A _10477_/B _10481_/A vssd1 vssd1 vccd1 vccd1 _15531_/D sky130_fd_sc_hd__nor3_1
X_15004_ _15001_/X _14996_/A _14999_/B _15003_/Y vssd1 vssd1 vccd1 vccd1 _16319_/D
+ sky130_fd_sc_hd__o31a_1
X_12216_ _15804_/Q _12270_/B _12216_/C vssd1 vssd1 vccd1 vccd1 _12216_/Y sky130_fd_sc_hd__nand3_1
X_13196_ _13202_/B _13196_/B vssd1 vssd1 vccd1 vccd1 _13198_/A sky130_fd_sc_hd__or2_1
X_12147_ _12147_/A _12147_/B _12147_/C vssd1 vssd1 vccd1 vccd1 _12148_/C sky130_fd_sc_hd__nand3_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12078_ _12092_/C vssd1 vssd1 vccd1 vccd1 _12102_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11029_ _11036_/B _11029_/B vssd1 vssd1 vccd1 vccd1 _11031_/A sky130_fd_sc_hd__or2_1
X_15906_ _15907_/CLK _15906_/D vssd1 vssd1 vccd1 vccd1 _15906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15837_ _07603_/A _15837_/D vssd1 vssd1 vccd1 vccd1 _15837_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15768_ _15794_/CLK _15768_/D vssd1 vssd1 vccd1 vccd1 _15768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14719_ _16259_/Q _14717_/C _14718_/X vssd1 vssd1 vccd1 vccd1 _14720_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15699_ _15763_/CLK _15699_/D vssd1 vssd1 vccd1 vccd1 _15699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08249_/A sky130_fd_sc_hd__or2_1
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_15 _11078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _13693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 _13919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08171_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07955_ _10812_/A _07922_/B _07954_/Y vssd1 vssd1 vccd1 vccd1 _07979_/A sky130_fd_sc_hd__o21ai_2
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07886_ _07886_/A _07886_/B vssd1 vssd1 vccd1 vccd1 _07887_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09625_ _09623_/Y _09619_/C _09621_/X _09622_/Y vssd1 vssd1 vccd1 vccd1 _09626_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_56_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09556_ _10134_/A vssd1 vssd1 vccd1 vccd1 _09784_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08507_ _08505_/Y _08497_/C _08500_/X _08502_/Y vssd1 vssd1 vccd1 vccd1 _08508_/C
+ sky130_fd_sc_hd__a211o_1
X_09487_ _09487_/A _09487_/B _09493_/A vssd1 vssd1 vccd1 vccd1 _15378_/D sky130_fd_sc_hd__nor3_1
XFILLER_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08438_ _08435_/Y _08437_/X _08335_/X vssd1 vssd1 vccd1 vccd1 _08438_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_137_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ _15211_/Q _08403_/B vssd1 vssd1 vccd1 vccd1 _08371_/B sky130_fd_sc_hd__and2_1
X_10400_ _11551_/A vssd1 vssd1 vccd1 vccd1 _10629_/A sky130_fd_sc_hd__clkbuf_2
X_11380_ _11378_/A _11378_/B _11379_/X vssd1 vssd1 vccd1 vccd1 _15672_/D sky130_fd_sc_hd__a21oi_1
XFILLER_109_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10331_ _15511_/Q _10512_/B _10331_/C vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__and3_1
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10262_ _15500_/Q _10268_/C _10030_/X vssd1 vssd1 vccd1 vccd1 _10262_/Y sky130_fd_sc_hd__a21oi_1
X_13050_ _13050_/A vssd1 vssd1 vccd1 vccd1 _15938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12001_ _12569_/A vssd1 vssd1 vccd1 vccd1 _12001_/X sky130_fd_sc_hd__clkbuf_2
X_10193_ _10191_/X _10192_/Y _10188_/B _10189_/C vssd1 vssd1 vccd1 vccd1 _10195_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_120_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13952_ _13952_/A _13952_/B vssd1 vssd1 vccd1 vccd1 _13952_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _15913_/Q _13066_/B _12908_/C vssd1 vssd1 vccd1 vccd1 _12903_/Y sky130_fd_sc_hd__nand3_1
X_13883_ _13883_/A vssd1 vssd1 vccd1 vccd1 _16082_/D sky130_fd_sc_hd__clkbuf_1
X_15622_ _15194_/Q _15622_/D vssd1 vssd1 vccd1 vccd1 _15622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12834_ _12832_/X _12833_/Y _12829_/B _12830_/C vssd1 vssd1 vccd1 vccd1 _12836_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15655_/CLK _15553_/D vssd1 vssd1 vccd1 vccd1 _15553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12765_ _12786_/C vssd1 vssd1 vccd1 vccd1 _12798_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _16210_/Q _14525_/C _14503_/X vssd1 vssd1 vccd1 vccd1 _14506_/B sky130_fd_sc_hd__a21oi_1
X_11716_ _11722_/A _11714_/Y _11715_/Y _11708_/C vssd1 vssd1 vccd1 vccd1 _11718_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15484_ _15484_/CLK _15484_/D vssd1 vssd1 vccd1 vccd1 _15484_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12919_/A _12699_/C vssd1 vssd1 vccd1 vccd1 _12696_/X sky130_fd_sc_hd__or2_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ _16194_/Q _14474_/B _14435_/C vssd1 vssd1 vccd1 vccd1 _14442_/A sky130_fd_sc_hd__and3_1
X_11647_ _11647_/A vssd1 vssd1 vccd1 vccd1 _15714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14366_ _14533_/A _14366_/B vssd1 vssd1 vccd1 vccd1 _14366_/Y sky130_fd_sc_hd__nor2_1
X_11578_ _11576_/X _11577_/Y _11573_/B _11574_/C vssd1 vssd1 vccd1 vccd1 _11580_/B
+ sky130_fd_sc_hd__o211ai_1
X_16105_ _16222_/CLK _16105_/D vssd1 vssd1 vccd1 vccd1 _16105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13317_ _14287_/A vssd1 vssd1 vccd1 vccd1 _13317_/X sky130_fd_sc_hd__clkbuf_4
X_10529_ _10549_/C vssd1 vssd1 vccd1 vccd1 _10561_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14297_ _14297_/A vssd1 vssd1 vccd1 vccd1 _16163_/D sky130_fd_sc_hd__clkbuf_1
X_16036_ _16050_/CLK _16036_/D vssd1 vssd1 vccd1 vccd1 _16036_/Q sky130_fd_sc_hd__dfxtp_2
X_13248_ _13255_/B _13248_/B vssd1 vssd1 vccd1 vccd1 _13252_/A sky130_fd_sc_hd__or2_1
XFILLER_124_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13179_ _14993_/A vssd1 vssd1 vccd1 vccd1 _13179_/X sky130_fd_sc_hd__buf_2
XFILLER_123_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07740_ _07740_/A _07740_/B vssd1 vssd1 vccd1 vccd1 _08136_/B sky130_fd_sc_hd__xor2_4
XFILLER_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07671_ _12616_/A vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__buf_2
X_09410_ _09699_/A vssd1 vssd1 vccd1 vccd1 _09644_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09341_ _13693_/A vssd1 vssd1 vccd1 vccd1 _09572_/B sky130_fd_sc_hd__buf_2
XFILLER_40_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09272_ _09270_/X _09271_/Y _09266_/B _09267_/C vssd1 vssd1 vccd1 vccd1 _09274_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_139_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08223_ _08080_/A _08080_/B _08222_/Y vssd1 vssd1 vccd1 vccd1 _08300_/B sky130_fd_sc_hd__a21o_2
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08154_ _08175_/A _08175_/B vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__xor2_4
XFILLER_107_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08085_ _13097_/C _07756_/B _07755_/A vssd1 vssd1 vccd1 vccd1 _08104_/A sky130_fd_sc_hd__o21ai_4
XFILLER_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08987_ _15302_/Q _09158_/B _08989_/C vssd1 vssd1 vccd1 vccd1 _08987_/X sky130_fd_sc_hd__and3_1
XFILLER_29_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07938_ _08731_/A _08160_/B vssd1 vssd1 vccd1 vccd1 _07939_/B sky130_fd_sc_hd__xnor2_2
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07869_ _12304_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _08016_/A sky130_fd_sc_hd__xnor2_2
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09608_ _09643_/A _09608_/B _09612_/A vssd1 vssd1 vccd1 vccd1 _15396_/D sky130_fd_sc_hd__nor3_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ _10902_/A _10880_/B _10880_/C vssd1 vssd1 vccd1 vccd1 _10881_/A sky130_fd_sc_hd__and3_1
XFILLER_43_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09539_ _09575_/A _09539_/B _09539_/C vssd1 vssd1 vccd1 vccd1 _09540_/A sky130_fd_sc_hd__and3_1
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ _12565_/A _12550_/B _12550_/C vssd1 vssd1 vccd1 vccd1 _12551_/A sky130_fd_sc_hd__and3_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _15700_/Q _15699_/Q _15698_/Q _11273_/X vssd1 vssd1 vccd1 vccd1 _15692_/D
+ sky130_fd_sc_hd__o31a_1
X_12481_ _13041_/A vssd1 vssd1 vccd1 vccd1 _12481_/X sky130_fd_sc_hd__buf_2
X_14220_ _14304_/A _14220_/B _14223_/B vssd1 vssd1 vccd1 vccd1 _16146_/D sky130_fd_sc_hd__nor3_1
X_11432_ _15682_/Q _11431_/C _11199_/X vssd1 vssd1 vccd1 vccd1 _11433_/B sky130_fd_sc_hd__a21oi_1
XFILLER_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _13920_/X _14146_/B _14150_/Y vssd1 vssd1 vccd1 vccd1 _16132_/D sky130_fd_sc_hd__o21a_1
X_11363_ _11360_/X _11361_/Y _11362_/Y _11358_/C vssd1 vssd1 vccd1 vccd1 _11365_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_138_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _13679_/A vssd1 vssd1 vccd1 vccd1 _14250_/A sky130_fd_sc_hd__buf_2
XFILLER_125_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10314_ _10312_/Y _10308_/C _10310_/X _10311_/Y vssd1 vssd1 vccd1 vccd1 _10315_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14082_ _14080_/X _14081_/Y _14077_/B _14078_/C vssd1 vssd1 vccd1 vccd1 _14084_/B
+ sky130_fd_sc_hd__o211ai_1
X_11294_ _11294_/A vssd1 vssd1 vccd1 vccd1 _15659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _13069_/A _13033_/B _13033_/C vssd1 vssd1 vccd1 vccd1 _13034_/A sky130_fd_sc_hd__and3_1
X_10245_ _10266_/A _10245_/B _10245_/C vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__and3_1
XFILLER_133_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10176_ _15493_/Q _15492_/Q _15491_/Q _10119_/X vssd1 vssd1 vccd1 vccd1 _15485_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14984_ _14984_/A _14984_/B _14984_/C vssd1 vssd1 vccd1 vccd1 _14985_/C sky130_fd_sc_hd__nand3_1
XFILLER_120_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13935_ _13945_/C vssd1 vssd1 vccd1 vccd1 _13957_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13866_ _13666_/X _13863_/C _13865_/Y vssd1 vssd1 vccd1 vccd1 _16079_/D sky130_fd_sc_hd__a21oi_1
X_15605_ _15194_/Q _15605_/D vssd1 vssd1 vccd1 vccd1 _15605_/Q sky130_fd_sc_hd__dfxtp_1
X_12817_ _15907_/Q _15906_/Q _15905_/Q _12704_/X vssd1 vssd1 vccd1 vccd1 _15899_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13797_ _13844_/A _13797_/B _13797_/C vssd1 vssd1 vccd1 vccd1 _13798_/A sky130_fd_sc_hd__and3_1
XFILLER_43_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15536_ _15655_/CLK _15536_/D vssd1 vssd1 vccd1 vccd1 _15536_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _15889_/Q _12861_/B _12748_/C vssd1 vssd1 vccd1 vccd1 _12757_/B sky130_fd_sc_hd__and3_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15467_ _15485_/CLK _15467_/D vssd1 vssd1 vccd1 vccd1 _15467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12679_ _12677_/Y _12673_/C _12675_/X _12676_/Y vssd1 vssd1 vccd1 vccd1 _12680_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14418_ _14325_/X _14411_/B _14326_/X vssd1 vssd1 vccd1 vccd1 _14420_/A sky130_fd_sc_hd__a21oi_1
X_15398_ _15483_/CLK _15398_/D vssd1 vssd1 vccd1 vccd1 _15398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14349_ _14427_/A _14349_/B _14352_/B vssd1 vssd1 vccd1 vccd1 _16173_/D sky130_fd_sc_hd__nor3_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16019_ _16031_/CLK _16019_/D vssd1 vssd1 vccd1 vccd1 _16019_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_143_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08910_ _10354_/A vssd1 vssd1 vccd1 vccd1 _10065_/A sky130_fd_sc_hd__buf_4
X_09890_ _09903_/C vssd1 vssd1 vccd1 vccd1 _09911_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08878_/A _08841_/B _08841_/C vssd1 vssd1 vccd1 vccd1 _08842_/A sky130_fd_sc_hd__and3_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08778_/A _08770_/Y _08771_/Y _08765_/C vssd1 vssd1 vccd1 vccd1 _08774_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07723_ _08127_/A _08128_/B vssd1 vssd1 vccd1 vccd1 _07729_/A sky130_fd_sc_hd__xnor2_4
XFILLER_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07654_ input4/X vssd1 vssd1 vccd1 vccd1 _12726_/A sky130_fd_sc_hd__buf_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ _09345_/A _09324_/B _09324_/C vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__and3_1
XFILLER_34_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09255_ _15359_/Q _15358_/Q _15357_/Q _09194_/X vssd1 vssd1 vccd1 vccd1 _15342_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_138_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08206_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08206_/X sky130_fd_sc_hd__and2_1
X_09186_ _09184_/A _09184_/B _09185_/X vssd1 vssd1 vccd1 vccd1 _15331_/D sky130_fd_sc_hd__a21oi_1
XFILLER_4_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08137_ _07757_/A _07757_/B _08136_/Y vssd1 vssd1 vccd1 vccd1 _08252_/B sky130_fd_sc_hd__o21a_2
XFILLER_107_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08068_ _07780_/A _07780_/B _07779_/A vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__o21ai_1
XFILLER_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10030_ _10610_/A vssd1 vssd1 vccd1 vccd1 _10030_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ _11975_/B _11976_/C _11978_/X _11979_/Y vssd1 vssd1 vccd1 vccd1 _11982_/C
+ sky130_fd_sc_hd__a211o_1
X_13720_ _13720_/A vssd1 vssd1 vccd1 vccd1 _13720_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10932_ _15605_/Q _10939_/B _13526_/A vssd1 vssd1 vccd1 vccd1 _10936_/B sky130_fd_sc_hd__nand3_1
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13651_ _13658_/A _13649_/Y _13650_/Y _13646_/C vssd1 vssd1 vccd1 vccd1 _13653_/B
+ sky130_fd_sc_hd__o211a_1
X_10863_ _10863_/A _10863_/B _10863_/C vssd1 vssd1 vccd1 vccd1 _10865_/B sky130_fd_sc_hd__or3_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12602_ _15867_/Q _12610_/C _12377_/X vssd1 vssd1 vccd1 vccd1 _12602_/Y sky130_fd_sc_hd__a21oi_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A vssd1 vssd1 vccd1 vccd1 _16028_/D sky130_fd_sc_hd__clkbuf_1
X_10794_ _15581_/Q _11023_/B _10798_/C vssd1 vssd1 vccd1 vccd1 _10794_/Y sky130_fd_sc_hd__nand3_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15339_/CLK _15321_/D vssd1 vssd1 vccd1 vccd1 _15321_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12533_ _15854_/Q vssd1 vssd1 vccd1 vccd1 _12546_/C sky130_fd_sc_hd__inv_2
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15252_ _15260_/CLK _15252_/D vssd1 vssd1 vccd1 vccd1 _15252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12464_ _12471_/B _12464_/B vssd1 vssd1 vccd1 vccd1 _12466_/A sky130_fd_sc_hd__or2_1
X_14203_ _16158_/Q _16160_/Q _16159_/Q _14202_/X vssd1 vssd1 vccd1 vccd1 _16143_/D
+ sky130_fd_sc_hd__o31a_1
X_11415_ _15680_/Q _11423_/C _11184_/X vssd1 vssd1 vccd1 vccd1 _11415_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_125_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15183_ _15178_/A _15181_/B _15043_/X vssd1 vssd1 vccd1 vccd1 _15189_/C sky130_fd_sc_hd__o21a_1
X_12395_ _12393_/Y _12389_/C _12391_/X _12392_/Y vssd1 vssd1 vccd1 vccd1 _12396_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14134_ _14133_/X _14132_/Y _14042_/X vssd1 vssd1 vccd1 vccd1 _14134_/Y sky130_fd_sc_hd__a21oi_1
X_11346_ _11634_/A vssd1 vssd1 vccd1 vccd1 _11576_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_140_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14065_ _16071_/Q vssd1 vssd1 vccd1 vccd1 _14071_/C sky130_fd_sc_hd__inv_2
XFILLER_125_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11277_ _11298_/C vssd1 vssd1 vccd1 vccd1 _11311_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13016_ _15933_/Q _13071_/B _13016_/C vssd1 vssd1 vccd1 vccd1 _13025_/A sky130_fd_sc_hd__and3_1
X_10228_ _10284_/A _10228_/B _10228_/C vssd1 vssd1 vccd1 vccd1 _10230_/B sky130_fd_sc_hd__or3_1
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10159_ _10165_/A _10156_/Y _10158_/Y _10153_/C vssd1 vssd1 vccd1 vccd1 _10161_/B
+ sky130_fd_sc_hd__o211a_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_14967_ _15051_/A _15010_/B _14967_/C vssd1 vssd1 vccd1 vccd1 _14969_/A sky130_fd_sc_hd__and3_1
X_13918_ _13912_/X _13916_/B _13917_/Y vssd1 vssd1 vccd1 vccd1 _16086_/D sky130_fd_sc_hd__o21a_1
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14898_ _16313_/Q _16312_/Q _16311_/Q _14818_/X vssd1 vssd1 vccd1 vccd1 _16296_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13849_ _16077_/Q _14095_/B _13853_/C vssd1 vssd1 vccd1 vccd1 _13849_/Y sky130_fd_sc_hd__nand3_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15519_ _15655_/CLK _15519_/D vssd1 vssd1 vccd1 vccd1 _15519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09040_ _15310_/Q _09047_/C _08920_/X vssd1 vssd1 vccd1 vccd1 _09040_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _09942_/A vssd1 vssd1 vccd1 vccd1 _15448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _09930_/A _09873_/B _09877_/B vssd1 vssd1 vccd1 vccd1 _15437_/D sky130_fd_sc_hd__nor3_1
XFILLER_58_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _09693_/A vssd1 vssd1 vccd1 vccd1 _08824_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08755_ _08753_/Y _08749_/C _08751_/X _08752_/Y vssd1 vssd1 vccd1 vccd1 _08756_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_66_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07706_ _14326_/A vssd1 vssd1 vccd1 vccd1 _14814_/A sky130_fd_sc_hd__buf_2
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08686_ _15256_/Q _08919_/B _08686_/C vssd1 vssd1 vccd1 vccd1 _08686_/X sky130_fd_sc_hd__and3_1
XFILLER_26_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _07638_/B _07638_/C _07638_/A vssd1 vssd1 vccd1 vccd1 _07639_/B sky130_fd_sc_hd__a21o_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09307_ _14372_/A vssd1 vssd1 vccd1 vccd1 _09307_/X sky130_fd_sc_hd__buf_2
XFILLER_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ _15339_/Q _09238_/B _09242_/C vssd1 vssd1 vccd1 vccd1 _09238_/Y sky130_fd_sc_hd__nand3_1
XFILLER_108_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09169_ _09165_/X _09167_/Y _09168_/Y _09163_/C vssd1 vssd1 vccd1 vccd1 _09171_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_107_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11200_ _15646_/Q _11198_/C _11199_/X vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__a21oi_1
XFILLER_135_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12180_ _12187_/B _12180_/B vssd1 vssd1 vccd1 vccd1 _12182_/A sky130_fd_sc_hd__or2_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11131_ _11126_/X _11127_/Y _11130_/Y _11124_/C vssd1 vssd1 vccd1 vccd1 _11133_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_134_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11062_ _11076_/A _11062_/B _11062_/C vssd1 vssd1 vccd1 vccd1 _11063_/A sky130_fd_sc_hd__and3_1
XFILLER_135_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10013_ _10013_/A _10013_/B _10013_/C vssd1 vssd1 vccd1 vccd1 _10014_/C sky130_fd_sc_hd__nand3_1
XFILLER_49_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15870_ _15907_/CLK _15870_/D vssd1 vssd1 vccd1 vccd1 _15870_/Q sky130_fd_sc_hd__dfxtp_1
X_14821_ _14826_/C vssd1 vssd1 vccd1 vccd1 _14838_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14752_ _14758_/A _14751_/Y _14747_/B _14748_/C vssd1 vssd1 vccd1 vccd1 _14754_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11964_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12084_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13703_ _16050_/Q _13801_/B _13707_/C vssd1 vssd1 vccd1 vccd1 _13703_/Y sky130_fd_sc_hd__nand3_1
X_10915_ _10915_/A _10915_/B vssd1 vssd1 vccd1 vccd1 _10920_/C sky130_fd_sc_hd__nor2_1
X_14683_ _14843_/A _14683_/B vssd1 vssd1 vccd1 vccd1 _14683_/X sky130_fd_sc_hd__or2_1
XFILLER_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11895_ _11895_/A _11895_/B vssd1 vssd1 vccd1 vccd1 _11901_/C sky130_fd_sc_hd__nor2_1
X_13634_ _16040_/Q _13738_/B _13634_/C vssd1 vssd1 vccd1 vccd1 _13634_/X sky130_fd_sc_hd__and3_1
XFILLER_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10846_ _10846_/A vssd1 vssd1 vccd1 vccd1 _15589_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16353_ _16353_/CLK _16353_/D vssd1 vssd1 vccd1 vccd1 _16353_/Q sky130_fd_sc_hd__dfxtp_2
X_13565_ _13565_/A vssd1 vssd1 vccd1 vccd1 _16024_/D sky130_fd_sc_hd__clkbuf_1
X_10777_ _15580_/Q _10778_/C _10663_/X vssd1 vssd1 vccd1 vccd1 _10777_/Y sky130_fd_sc_hd__a21oi_1
X_15304_ _15322_/CLK _15304_/D vssd1 vssd1 vccd1 vccd1 _15304_/Q sky130_fd_sc_hd__dfxtp_1
X_12516_ _12522_/A _12513_/Y _12515_/Y _12510_/C vssd1 vssd1 vccd1 vccd1 _12518_/B
+ sky130_fd_sc_hd__o211a_1
X_16284_ _16321_/CLK _16284_/D vssd1 vssd1 vccd1 vccd1 _16284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13496_ _13496_/A vssd1 vssd1 vccd1 vccd1 _16012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15235_ _15351_/CLK _15235_/D vssd1 vssd1 vccd1 vccd1 _15235_/Q sky130_fd_sc_hd__dfxtp_2
X_12447_ _12447_/A vssd1 vssd1 vccd1 vccd1 _15840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15166_ _16365_/Q _15165_/C _13981_/B vssd1 vssd1 vccd1 vccd1 _15168_/C sky130_fd_sc_hd__a21o_1
X_12378_ _15831_/Q _12386_/C _12377_/X vssd1 vssd1 vccd1 vccd1 _12378_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_125_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14117_ _16129_/Q _14117_/B _14117_/C vssd1 vssd1 vccd1 vccd1 _14122_/A sky130_fd_sc_hd__and3_1
XFILLER_126_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11329_ _11365_/A _11329_/B _11329_/C vssd1 vssd1 vccd1 vccd1 _11330_/A sky130_fd_sc_hd__and3_1
X_15097_ _16347_/Q _15096_/C _14942_/X vssd1 vssd1 vccd1 vccd1 _15099_/C sky130_fd_sc_hd__a21o_1
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14048_ _14046_/X _14048_/B vssd1 vssd1 vccd1 vccd1 _14048_/X sky130_fd_sc_hd__and2b_1
XFILLER_95_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15999_ _16022_/CLK _15999_/D vssd1 vssd1 vccd1 vccd1 _15999_/Q sky130_fd_sc_hd__dfxtp_2
X_08540_ _12758_/A _08540_/B _08540_/C vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__or3_1
XFILLER_63_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08471_ _15224_/Q _08471_/B vssd1 vssd1 vccd1 vccd1 _15224_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09023_ _15323_/Q _15322_/Q _15321_/Q _08901_/X vssd1 vssd1 vccd1 vccd1 _15306_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_136_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09925_ _15447_/Q _10155_/B _09925_/C vssd1 vssd1 vccd1 vccd1 _09934_/A sky130_fd_sc_hd__and3_1
XFILLER_120_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09856_ _09853_/X _09854_/Y _09855_/Y _09851_/C vssd1 vssd1 vccd1 vccd1 _09858_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _08807_/A vssd1 vssd1 vccd1 vccd1 _15273_/D sky130_fd_sc_hd__clkbuf_1
X_09787_ _15426_/Q _09796_/C _09786_/X vssd1 vssd1 vccd1 vccd1 _09787_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _08774_/A _08738_/B _08742_/A vssd1 vssd1 vccd1 vccd1 _15262_/D sky130_fd_sc_hd__nor3_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _08704_/A _08669_/B _08669_/C vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__and3_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10700_/A vssd1 vssd1 vccd1 vccd1 _10714_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _15721_/Q _11719_/C _11624_/X vssd1 vssd1 vccd1 vccd1 _11682_/B sky130_fd_sc_hd__a21oi_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _10693_/A vssd1 vssd1 vccd1 vccd1 _10676_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13350_ _15989_/Q _13349_/C _13194_/X vssd1 vssd1 vccd1 vccd1 _13351_/B sky130_fd_sc_hd__a21oi_1
XFILLER_139_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10562_ _11137_/A vssd1 vssd1 vccd1 vccd1 _10562_/X sky130_fd_sc_hd__buf_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _12337_/A _12301_/B _12301_/C vssd1 vssd1 vccd1 vccd1 _12302_/A sky130_fd_sc_hd__and3_1
X_13281_ _13281_/A _13281_/B _13281_/C vssd1 vssd1 vccd1 vccd1 _13282_/A sky130_fd_sc_hd__and3_1
XFILLER_139_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10493_ _10490_/X _10491_/Y _10492_/Y _10488_/C vssd1 vssd1 vccd1 vccd1 _10495_/B
+ sky130_fd_sc_hd__o211ai_1
X_15020_ _16328_/Q _15036_/C _14901_/X vssd1 vssd1 vccd1 vccd1 _15023_/B sky130_fd_sc_hd__a21oi_1
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12232_ _12238_/A _12229_/Y _12231_/Y _12226_/C vssd1 vssd1 vccd1 vccd1 _12234_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _12163_/A vssd1 vssd1 vccd1 vccd1 _15795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11114_ _15633_/Q _11121_/C _10940_/X vssd1 vssd1 vccd1 vccd1 _11114_/Y sky130_fd_sc_hd__a21oi_1
X_12094_ _15786_/Q _12102_/C _12093_/X vssd1 vssd1 vccd1 vccd1 _12094_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11045_ _11066_/C vssd1 vssd1 vccd1 vccd1 _11078_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15922_ _07603_/A _15922_/D vssd1 vssd1 vccd1 vccd1 _15922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ _15907_/CLK _15853_/D vssd1 vssd1 vccd1 vccd1 _15853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14804_ _14847_/A _14811_/C vssd1 vssd1 vccd1 vccd1 _14804_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12996_ _15930_/Q _12996_/B _12996_/C vssd1 vssd1 vccd1 vccd1 _12996_/X sky130_fd_sc_hd__and3_1
X_15784_ _15794_/CLK _15784_/D vssd1 vssd1 vccd1 vccd1 _15784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11947_ _11953_/A _11944_/Y _11946_/Y _11941_/C vssd1 vssd1 vccd1 vccd1 _11949_/B
+ sky130_fd_sc_hd__o211a_1
X_14735_ _07707_/X _14733_/A _14734_/Y vssd1 vssd1 vccd1 vccd1 _16259_/D sky130_fd_sc_hd__o21a_1
XFILLER_45_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14666_ _16248_/Q _14665_/C _15165_/B vssd1 vssd1 vccd1 vccd1 _14668_/C sky130_fd_sc_hd__a21o_1
X_11878_ _15752_/Q _12107_/B _11885_/C vssd1 vssd1 vccd1 vccd1 _11878_/X sky130_fd_sc_hd__and3_1
X_13617_ _13617_/A vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__clkbuf_2
X_10829_ _10845_/A _10829_/B _10829_/C vssd1 vssd1 vccd1 vccd1 _10830_/A sky130_fd_sc_hd__and3_1
X_14597_ _14626_/A _14597_/B _14600_/B vssd1 vssd1 vccd1 vccd1 _16227_/D sky130_fd_sc_hd__nor3_1
XFILLER_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16336_ _16337_/CLK _16336_/D vssd1 vssd1 vccd1 vccd1 _16336_/Q sky130_fd_sc_hd__dfxtp_2
X_13548_ _16024_/Q _13648_/B _13548_/C vssd1 vssd1 vccd1 vccd1 _13557_/A sky130_fd_sc_hd__and3_1
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16267_ _16268_/CLK _16267_/D vssd1 vssd1 vccd1 vccd1 _16267_/Q sky130_fd_sc_hd__dfxtp_1
X_13479_ _13480_/B _13480_/C _13480_/A vssd1 vssd1 vccd1 vccd1 _13481_/B sky130_fd_sc_hd__a21o_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15218_ _16224_/CLK _15218_/D vssd1 vssd1 vccd1 vccd1 state1[3] sky130_fd_sc_hd__dfxtp_2
X_16198_ _16247_/CLK _16198_/D vssd1 vssd1 vccd1 vccd1 _16198_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _15144_/A _15147_/B _15043_/X vssd1 vssd1 vccd1 vccd1 _15155_/C sky130_fd_sc_hd__o21a_1
XFILLER_114_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ _07909_/A _07909_/B _07970_/X vssd1 vssd1 vccd1 vccd1 _07973_/B sky130_fd_sc_hd__o21a_1
XFILLER_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09710_ _09746_/A _09710_/B _09710_/C vssd1 vssd1 vccd1 vccd1 _09711_/A sky130_fd_sc_hd__and3_1
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09641_ _09647_/A _09639_/Y _09640_/Y _09635_/C vssd1 vssd1 vccd1 vccd1 _09643_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09572_ _15391_/Q _09572_/B _09577_/C vssd1 vssd1 vccd1 vccd1 _09572_/Y sky130_fd_sc_hd__nand3_1
XFILLER_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08523_ _11424_/A vssd1 vssd1 vccd1 vccd1 _09693_/A sky130_fd_sc_hd__buf_2
XFILLER_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08454_ _08443_/A _08448_/A _08465_/A _08453_/Y vssd1 vssd1 vccd1 vccd1 _08456_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08385_ _08386_/B _08386_/C _08386_/A vssd1 vssd1 vccd1 vccd1 _08387_/A sky130_fd_sc_hd__a21oi_1
XFILLER_149_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09006_ _09004_/Y _08999_/C _09011_/A _09002_/Y vssd1 vssd1 vccd1 vccd1 _09011_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_136_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09908_ _09908_/A vssd1 vssd1 vccd1 vccd1 _15443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09839_ _09930_/A _09839_/B _09843_/A vssd1 vssd1 vccd1 vccd1 _15432_/D sky130_fd_sc_hd__nor3_1
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12850_ _12848_/Y _12843_/C _12845_/X _12846_/Y vssd1 vssd1 vccd1 vccd1 _12851_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _11801_/A _11801_/B _11801_/C vssd1 vssd1 vccd1 vccd1 _11802_/C sky130_fd_sc_hd__nand3_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12781_ _12774_/B _12775_/C _12778_/X _12779_/Y vssd1 vssd1 vccd1 vccd1 _12782_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14520_/A _14520_/B vssd1 vssd1 vccd1 vccd1 _14520_/Y sky130_fd_sc_hd__nor2_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ _15728_/Q vssd1 vssd1 vccd1 vccd1 _11745_/C sky130_fd_sc_hd__inv_2
XFILLER_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14446_/Y _14449_/X _14450_/Y vssd1 vssd1 vccd1 vccd1 _16193_/D sky130_fd_sc_hd__o21a_1
X_11663_ _15718_/Q _11662_/C _11488_/X vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__a21oi_1
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _15998_/Q _13401_/C _13194_/X vssd1 vssd1 vccd1 vccd1 _13403_/B sky130_fd_sc_hd__a21oi_1
X_10614_ _10612_/Y _10607_/C _10609_/X _10611_/Y vssd1 vssd1 vccd1 vccd1 _10615_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14382_ _14979_/A vssd1 vssd1 vccd1 vccd1 _14552_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11594_ _15706_/Q _11650_/B _11599_/C vssd1 vssd1 vccd1 vccd1 _11594_/Y sky130_fd_sc_hd__nand3_1
X_16121_ _16123_/CLK _16121_/D vssd1 vssd1 vccd1 vccd1 _16121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13333_ _15987_/Q _13333_/B _13341_/C vssd1 vssd1 vccd1 vccd1 _13333_/X sky130_fd_sc_hd__and3_1
XFILLER_127_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ _10545_/A vssd1 vssd1 vccd1 vccd1 _15542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16052_ _16052_/CLK _16052_/D vssd1 vssd1 vccd1 vccd1 _16052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13264_ _13291_/C vssd1 vssd1 vccd1 vccd1 _13297_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10476_ _15532_/Q _10532_/B _10484_/C vssd1 vssd1 vccd1 vccd1 _10481_/A sky130_fd_sc_hd__and3_1
X_15003_ _15045_/A _15010_/C vssd1 vssd1 vccd1 vccd1 _15003_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12215_ _15805_/Q _12216_/C _12100_/X vssd1 vssd1 vccd1 vccd1 _12215_/Y sky130_fd_sc_hd__a21oi_1
X_13195_ _15962_/Q _13193_/C _13194_/X vssd1 vssd1 vccd1 vccd1 _13196_/B sky130_fd_sc_hd__a21oi_1
XFILLER_123_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12146_ _12147_/B _12147_/C _12147_/A vssd1 vssd1 vccd1 vccd1 _12148_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ _12077_/A vssd1 vssd1 vccd1 vccd1 _12092_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11028_ _15619_/Q _11027_/C _10911_/X vssd1 vssd1 vccd1 vccd1 _11029_/B sky130_fd_sc_hd__a21oi_1
X_15905_ _15907_/CLK _15905_/D vssd1 vssd1 vccd1 vccd1 _15905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15836_ _15845_/CLK _15836_/D vssd1 vssd1 vccd1 vccd1 _15836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15767_ _15794_/CLK _15767_/D vssd1 vssd1 vccd1 vccd1 _15767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12979_ _13014_/A _12979_/B _12979_/C vssd1 vssd1 vccd1 vccd1 _12980_/A sky130_fd_sc_hd__and3_1
X_14718_ _15176_/B vssd1 vssd1 vccd1 vccd1 _14718_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15698_ _15794_/CLK _15698_/D vssd1 vssd1 vccd1 vccd1 _15698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14649_ _07675_/X _14641_/A _14644_/B _14648_/Y vssd1 vssd1 vccd1 vccd1 _16238_/D
+ sky130_fd_sc_hd__o31a_1
XANTENNA_16 _14869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_27 _11963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _14466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _07946_/C _08166_/Y _08169_/Y vssd1 vssd1 vccd1 vccd1 _15207_/D sky130_fd_sc_hd__o21a_1
XFILLER_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16319_ _16327_/CLK _16319_/D vssd1 vssd1 vccd1 vccd1 _16319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07954_ _15602_/Q _07954_/B vssd1 vssd1 vccd1 vccd1 _07954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07885_ _15620_/Q _07885_/B vssd1 vssd1 vccd1 vccd1 _07886_/B sky130_fd_sc_hd__or2_1
XFILLER_28_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09624_ _09621_/X _09622_/Y _09623_/Y _09619_/C vssd1 vssd1 vccd1 vccd1 _09626_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ _09555_/A vssd1 vssd1 vccd1 vccd1 _15388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08506_ _08500_/X _08502_/Y _08505_/Y _08497_/C vssd1 vssd1 vccd1 vccd1 _08508_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ _15379_/Q _09663_/B _09496_/C vssd1 vssd1 vccd1 vccd1 _09493_/A sky130_fd_sc_hd__and3_1
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08437_ _08428_/Y _08430_/Y _08436_/Y vssd1 vssd1 vccd1 vccd1 _08437_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08368_ _08368_/A _08368_/B vssd1 vssd1 vccd1 vccd1 _08442_/A sky130_fd_sc_hd__xor2_2
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08299_ _08219_/A _08219_/B _08218_/A vssd1 vssd1 vccd1 vccd1 _08304_/A sky130_fd_sc_hd__a21o_1
XFILLER_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10330_ _10353_/A _10330_/B _10336_/B vssd1 vssd1 vccd1 vccd1 _15509_/D sky130_fd_sc_hd__nor3_1
X_10261_ _15500_/Q _10317_/B _10268_/C vssd1 vssd1 vccd1 vccd1 _10261_/X sky130_fd_sc_hd__and3_1
XFILLER_127_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12000_ _15771_/Q _12228_/B _12000_/C vssd1 vssd1 vccd1 vccd1 _12010_/A sky130_fd_sc_hd__and3_1
XFILLER_133_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10192_ _15489_/Q _10199_/C _10075_/X vssd1 vssd1 vccd1 vccd1 _10192_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13951_ _16096_/Q _13957_/C _13893_/X vssd1 vssd1 vccd1 vccd1 _13953_/B sky130_fd_sc_hd__a21oi_1
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12902_ _15914_/Q _12908_/C _07672_/A vssd1 vssd1 vccd1 vccd1 _12902_/Y sky130_fd_sc_hd__a21oi_1
X_13882_ _14029_/A _13882_/B _13882_/C vssd1 vssd1 vccd1 vccd1 _13883_/A sky130_fd_sc_hd__and3_1
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15621_ _15194_/Q _15621_/D vssd1 vssd1 vccd1 vccd1 _15621_/Q sky130_fd_sc_hd__dfxtp_2
X_12833_ _15903_/Q _12840_/C _12661_/X vssd1 vssd1 vccd1 vccd1 _12833_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15655_/CLK _15552_/D vssd1 vssd1 vccd1 vccd1 _15552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12778_/C vssd1 vssd1 vccd1 vccd1 _12786_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11715_ _15725_/Q _11887_/B _11719_/C vssd1 vssd1 vccd1 vccd1 _11715_/Y sky130_fd_sc_hd__nand3_1
X_14503_ _14901_/A vssd1 vssd1 vccd1 vccd1 _14503_/X sky130_fd_sc_hd__buf_2
X_15483_ _15483_/CLK _15483_/D vssd1 vssd1 vccd1 vccd1 _15483_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12695_/A _12695_/B vssd1 vssd1 vccd1 vccd1 _12699_/C sky130_fd_sc_hd__nor2_1
XFILLER_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11646_ _11653_/A _11646_/B _11646_/C vssd1 vssd1 vccd1 vccd1 _11647_/A sky130_fd_sc_hd__and3_1
X_14434_ _14434_/A vssd1 vssd1 vccd1 vccd1 _14517_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14365_ _14532_/A _14365_/B vssd1 vssd1 vccd1 vccd1 _14366_/B sky130_fd_sc_hd__and2_1
X_11577_ _15705_/Q _11585_/C _11519_/X vssd1 vssd1 vccd1 vccd1 _11577_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13316_ _13316_/A vssd1 vssd1 vccd1 vccd1 _14287_/A sky130_fd_sc_hd__buf_4
X_16104_ _16114_/CLK _16104_/D vssd1 vssd1 vccd1 vccd1 _16104_/Q sky130_fd_sc_hd__dfxtp_1
X_10528_ _10540_/C vssd1 vssd1 vccd1 vccd1 _10549_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14296_ _14343_/A _14296_/B _14296_/C vssd1 vssd1 vccd1 vccd1 _14297_/A sky130_fd_sc_hd__and3_1
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13247_ _15971_/Q _13246_/C _13194_/X vssd1 vssd1 vccd1 vccd1 _13248_/B sky130_fd_sc_hd__a21oi_1
XFILLER_115_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16035_ _16060_/CLK _16035_/D vssd1 vssd1 vccd1 vccd1 _16035_/Q sky130_fd_sc_hd__dfxtp_1
X_10459_ _10457_/A _10457_/B _10458_/X vssd1 vssd1 vccd1 vccd1 _15528_/D sky130_fd_sc_hd__a21oi_1
XFILLER_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13178_ _15960_/Q _13333_/B _13187_/C vssd1 vssd1 vccd1 vccd1 _13178_/X sky130_fd_sc_hd__and3_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12129_ _12129_/A vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07670_ input5/X vssd1 vssd1 vccd1 vccd1 _12616_/A sky130_fd_sc_hd__buf_4
XFILLER_53_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15819_ _07603_/A _15819_/D vssd1 vssd1 vccd1 vccd1 _15819_/Q sky130_fd_sc_hd__dfxtp_2
X_09340_ _15357_/Q _09348_/C _09166_/X vssd1 vssd1 vccd1 vccd1 _09340_/Y sky130_fd_sc_hd__a21oi_1
X_09271_ _15346_/Q _09278_/C _09212_/X vssd1 vssd1 vccd1 vccd1 _09271_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08222_ _08222_/A _08222_/B vssd1 vssd1 vccd1 vccd1 _08222_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08153_ _07935_/A _07935_/B _08152_/Y vssd1 vssd1 vccd1 vccd1 _08175_/B sky130_fd_sc_hd__o21a_1
XFILLER_147_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08084_ _12983_/A _07767_/B _08083_/X vssd1 vssd1 vccd1 vccd1 _08105_/A sky130_fd_sc_hd__o21ai_4
XFILLER_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08986_ _08986_/A vssd1 vssd1 vccd1 vccd1 _15300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07937_ _08966_/A _07937_/B vssd1 vssd1 vccd1 vccd1 _08160_/B sky130_fd_sc_hd__xnor2_2
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07868_ _14022_/C _07868_/B vssd1 vssd1 vccd1 vccd1 _07869_/B sky130_fd_sc_hd__xnor2_2
XFILLER_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09607_ _15397_/Q _09663_/B _09615_/C vssd1 vssd1 vccd1 vccd1 _09612_/A sky130_fd_sc_hd__and3_1
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07799_ _12763_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _07800_/B sky130_fd_sc_hd__xnor2_2
X_09538_ _09537_/B _09537_/C _09307_/X vssd1 vssd1 vccd1 vccd1 _09539_/C sky130_fd_sc_hd__o21ai_1
X_09469_ _09476_/B _09469_/B vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__or2_1
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11500_ _11500_/A vssd1 vssd1 vccd1 vccd1 _15691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12480_ _12512_/C vssd1 vssd1 vccd1 vccd1 _12519_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _15682_/Q _11431_/B _11431_/C vssd1 vssd1 vccd1 vccd1 _11439_/B sky130_fd_sc_hd__and3_1
XFILLER_137_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14150_ _14149_/X _14146_/B _14049_/X vssd1 vssd1 vccd1 vccd1 _14150_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11362_ _15670_/Q _11362_/B _11367_/C vssd1 vssd1 vccd1 vccd1 _11362_/Y sky130_fd_sc_hd__nand3_1
X_13101_ _15949_/Q _14291_/A _13109_/C vssd1 vssd1 vccd1 vccd1 _13105_/B sky130_fd_sc_hd__nand3_1
X_10313_ _10310_/X _10311_/Y _10312_/Y _10308_/C vssd1 vssd1 vccd1 vccd1 _10315_/B
+ sky130_fd_sc_hd__o211ai_1
X_14081_ _16121_/Q _14080_/C _10950_/C vssd1 vssd1 vccd1 vccd1 _14081_/Y sky130_fd_sc_hd__a21oi_1
X_11293_ _11309_/A _11293_/B _11293_/C vssd1 vssd1 vccd1 vccd1 _11294_/A sky130_fd_sc_hd__and3_1
XFILLER_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _13031_/B _13031_/C _14970_/A vssd1 vssd1 vccd1 vccd1 _13033_/C sky130_fd_sc_hd__o21ai_1
X_10244_ _10244_/A _10244_/B _10244_/C vssd1 vssd1 vccd1 vccd1 _10245_/C sky130_fd_sc_hd__nand3_1
XFILLER_98_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10175_ _10175_/A vssd1 vssd1 vccd1 vccd1 _15484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14983_ _14984_/B _14984_/C _14984_/A vssd1 vssd1 vccd1 vccd1 _14985_/B sky130_fd_sc_hd__a21o_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13934_ _13937_/C vssd1 vssd1 vccd1 vccd1 _13945_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ _13666_/A _13863_/C _13720_/X vssd1 vssd1 vccd1 vccd1 _13865_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15604_ _15194_/Q _15604_/D vssd1 vssd1 vccd1 vccd1 _15604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12816_ _12816_/A vssd1 vssd1 vccd1 vccd1 _15898_/D sky130_fd_sc_hd__clkbuf_1
X_13796_ _13794_/Y _13789_/C _13792_/X _13793_/Y vssd1 vssd1 vccd1 vccd1 _13797_/C
+ sky130_fd_sc_hd__a211o_1
X_15535_ _15655_/CLK _15535_/D vssd1 vssd1 vccd1 vccd1 _15535_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12804_/A _12747_/B _12751_/B vssd1 vssd1 vccd1 vccd1 _15887_/D sky130_fd_sc_hd__nor3_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15466_ _15484_/CLK _15466_/D vssd1 vssd1 vccd1 vccd1 _15466_/Q sky130_fd_sc_hd__dfxtp_1
X_12678_ _12675_/X _12676_/Y _12677_/Y _12673_/C vssd1 vssd1 vccd1 vccd1 _12680_/B
+ sky130_fd_sc_hd__o211ai_1
X_11629_ _15713_/Q _11635_/C _11512_/X vssd1 vssd1 vccd1 vccd1 _11631_/C sky130_fd_sc_hd__a21o_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14417_ _14413_/X _14411_/B _14416_/Y vssd1 vssd1 vccd1 vccd1 _16186_/D sky130_fd_sc_hd__o21a_1
X_15397_ _15483_/CLK _15397_/D vssd1 vssd1 vccd1 vccd1 _15397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14348_ _14342_/B _14343_/C _14352_/A _14346_/Y vssd1 vssd1 vccd1 vccd1 _14352_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_6_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14279_ _14149_/X _14277_/B _14196_/X vssd1 vssd1 vccd1 vccd1 _14279_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16018_ _16022_/CLK _16018_/D vssd1 vssd1 vccd1 vccd1 _16018_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08839_/B _08839_/C _08726_/X vssd1 vssd1 vccd1 vccd1 _08841_/C sky130_fd_sc_hd__o21ai_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _15267_/Q _08947_/B _08775_/C vssd1 vssd1 vccd1 vccd1 _08771_/Y sky130_fd_sc_hd__nand3_1
XFILLER_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07722_ _15243_/Q _08125_/B vssd1 vssd1 vccd1 vccd1 _08128_/B sky130_fd_sc_hd__xnor2_2
XFILLER_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07653_ _08421_/A _07653_/B _07666_/B vssd1 vssd1 vccd1 vccd1 _15200_/D sky130_fd_sc_hd__nor3_1
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09323_ _09323_/A _09323_/B _09323_/C vssd1 vssd1 vccd1 vccd1 _09324_/C sky130_fd_sc_hd__nand3_1
XFILLER_80_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09254_ _09254_/A vssd1 vssd1 vccd1 vccd1 _15341_/D sky130_fd_sc_hd__clkbuf_1
X_08205_ _08205_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__nor2_1
X_09185_ _09185_/A _09190_/C vssd1 vssd1 vccd1 vccd1 _09185_/X sky130_fd_sc_hd__or2_1
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08136_ _15728_/Q _08136_/B vssd1 vssd1 vccd1 vccd1 _08136_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08067_ _14546_/C _07797_/B _08066_/X vssd1 vssd1 vccd1 vccd1 _08227_/B sky130_fd_sc_hd__o21ai_4
XFILLER_134_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08969_ _09001_/C vssd1 vssd1 vccd1 vccd1 _09008_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11980_ _11978_/X _11979_/Y _11975_/B _11976_/C vssd1 vssd1 vccd1 vccd1 _11982_/B
+ sky130_fd_sc_hd__o211ai_1
X_10931_ _10931_/A _10931_/B _10936_/A vssd1 vssd1 vccd1 vccd1 _15603_/D sky130_fd_sc_hd__nor3_1
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10862_ _10978_/A vssd1 vssd1 vccd1 vccd1 _10902_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13650_ _16041_/Q _13801_/B _13655_/C vssd1 vssd1 vccd1 vccd1 _13650_/Y sky130_fd_sc_hd__nand3_1
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12601_ _15867_/Q _12720_/B _12601_/C vssd1 vssd1 vccd1 vccd1 _12601_/X sky130_fd_sc_hd__and3_1
X_13581_ _13595_/A _13581_/B _13581_/C vssd1 vssd1 vccd1 vccd1 _13582_/A sky130_fd_sc_hd__and3_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _15582_/Q _10798_/C _10562_/X vssd1 vssd1 vccd1 vccd1 _10793_/Y sky130_fd_sc_hd__a21oi_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15320_ _15333_/CLK _15320_/D vssd1 vssd1 vccd1 vccd1 _15320_/Q sky130_fd_sc_hd__dfxtp_1
X_12532_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12652_/A sky130_fd_sc_hd__buf_2
XFILLER_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15251_ _15259_/CLK _15251_/D vssd1 vssd1 vccd1 vccd1 _15251_/Q sky130_fd_sc_hd__dfxtp_1
X_12463_ _15844_/Q _12462_/C _12347_/X vssd1 vssd1 vccd1 vccd1 _12464_/B sky130_fd_sc_hd__a21oi_1
XFILLER_138_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11414_ _15680_/Q _11533_/B _11423_/C vssd1 vssd1 vccd1 vccd1 _11414_/X sky130_fd_sc_hd__and3_1
X_14202_ _14818_/A vssd1 vssd1 vccd1 vccd1 _14202_/X sky130_fd_sc_hd__buf_2
X_15182_ _15180_/A _15180_/B _15181_/X vssd1 vssd1 vccd1 vccd1 _16363_/D sky130_fd_sc_hd__a21oi_1
X_12394_ _12391_/X _12392_/Y _12393_/Y _12389_/C vssd1 vssd1 vccd1 vccd1 _12396_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_125_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14133_ _14133_/A _14133_/B vssd1 vssd1 vccd1 vccd1 _14133_/X sky130_fd_sc_hd__or2_1
X_11345_ _11345_/A vssd1 vssd1 vccd1 vccd1 _15667_/D sky130_fd_sc_hd__clkbuf_1
X_14064_ _16133_/Q _16132_/Q _16131_/Q _13973_/X vssd1 vssd1 vccd1 vccd1 _16116_/D
+ sky130_fd_sc_hd__o31a_1
X_11276_ _11289_/C vssd1 vssd1 vccd1 vccd1 _11298_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13015_ _13015_/A vssd1 vssd1 vccd1 vccd1 _15931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10227_ _10404_/A vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10158_ _15482_/Q _10391_/B _10162_/C vssd1 vssd1 vccd1 vccd1 _10158_/Y sky130_fd_sc_hd__nand3_1
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_10089_ _10089_/A vssd1 vssd1 vccd1 vccd1 _15471_/D sky130_fd_sc_hd__clkbuf_1
X_14966_ _14966_/A _14966_/B vssd1 vssd1 vccd1 vccd1 _16311_/D sky130_fd_sc_hd__nor2_1
XFILLER_48_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13917_ _14054_/A _13917_/B vssd1 vssd1 vccd1 vccd1 _13917_/Y sky130_fd_sc_hd__nor2_1
X_14897_ _14814_/X _14895_/A _14896_/Y vssd1 vssd1 vccd1 vccd1 _16295_/D sky130_fd_sc_hd__o21a_1
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13848_ _16078_/Q _13853_/C _14270_/A vssd1 vssd1 vccd1 vccd1 _13848_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13779_ _16066_/Q _14074_/B _13785_/C vssd1 vssd1 vccd1 vccd1 _13782_/B sky130_fd_sc_hd__nand3_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15518_ _15655_/CLK _15518_/D vssd1 vssd1 vccd1 vccd1 _15518_/Q sky130_fd_sc_hd__dfxtp_1
X_15449_ _15449_/CLK _15449_/D vssd1 vssd1 vccd1 vccd1 _15449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09941_ _09977_/A _09941_/B _09941_/C vssd1 vssd1 vccd1 vccd1 _09942_/A sky130_fd_sc_hd__and3_1
XFILLER_131_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _09870_/Y _09865_/C _09877_/A _09868_/Y vssd1 vssd1 vccd1 vccd1 _09877_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08823_ _15277_/Q _09001_/B _08823_/C vssd1 vssd1 vccd1 vccd1 _08834_/A sky130_fd_sc_hd__and3_1
XFILLER_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08754_ _08751_/X _08752_/Y _08753_/Y _08749_/C vssd1 vssd1 vccd1 vccd1 _08756_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _12639_/A vssd1 vssd1 vccd1 vccd1 _14326_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _12661_/A vssd1 vssd1 vccd1 vccd1 _08919_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_92_clk _15584_/CLK vssd1 vssd1 vccd1 vccd1 _15575_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _15203_/Q _07633_/C _15165_/B vssd1 vssd1 vccd1 vccd1 _07638_/C sky130_fd_sc_hd__a21o_1
XFILLER_14_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09306_ _09419_/A _09306_/B _09306_/C vssd1 vssd1 vccd1 vccd1 _09309_/B sky130_fd_sc_hd__or3_1
XFILLER_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _15340_/Q _09242_/C _09118_/X vssd1 vssd1 vccd1 vccd1 _09237_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09168_ _15329_/Q _09285_/B _09173_/C vssd1 vssd1 vccd1 vccd1 _09168_/Y sky130_fd_sc_hd__nand3_1
XFILLER_108_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08119_ _15315_/Q vssd1 vssd1 vccd1 vccd1 _09138_/A sky130_fd_sc_hd__inv_2
XFILLER_119_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09099_ _09093_/B _09094_/C _09096_/X _09097_/Y vssd1 vssd1 vccd1 vccd1 _09100_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11130_ _15634_/Q _11362_/B _11136_/C vssd1 vssd1 vccd1 vccd1 _11130_/Y sky130_fd_sc_hd__nand3_1
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ _11054_/B _11055_/C _11058_/X _11059_/Y vssd1 vssd1 vccd1 vccd1 _11062_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_89_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10012_ _10013_/B _10013_/C _10013_/A vssd1 vssd1 vccd1 vccd1 _10014_/B sky130_fd_sc_hd__a21o_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14820_ _16269_/Q vssd1 vssd1 vccd1 vccd1 _14826_/C sky130_fd_sc_hd__inv_2
XFILLER_64_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14751_ _16267_/Q _14755_/C _07649_/X vssd1 vssd1 vccd1 vccd1 _14751_/Y sky130_fd_sc_hd__a21oi_1
X_11963_ _11963_/A vssd1 vssd1 vccd1 vccd1 _12532_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_83_clk clkbuf_opt_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15512_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13702_ _16051_/Q _13707_/C _13598_/X vssd1 vssd1 vccd1 vccd1 _13702_/Y sky130_fd_sc_hd__a21oi_1
X_10914_ _10914_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10915_/B sky130_fd_sc_hd__nor2_1
X_11894_ _11894_/A _11894_/B vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__nor2_1
X_14682_ _14682_/A _14682_/B vssd1 vssd1 vccd1 vccd1 _14683_/B sky130_fd_sc_hd__nor2_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13633_ _13633_/A vssd1 vssd1 vccd1 vccd1 _16037_/D sky130_fd_sc_hd__clkbuf_1
X_10845_ _10845_/A _10845_/B _10845_/C vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__and3_1
XFILLER_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16352_ _16352_/CLK _16352_/D vssd1 vssd1 vccd1 vccd1 _16352_/Q sky130_fd_sc_hd__dfxtp_2
X_10776_ _15580_/Q _10888_/B _10778_/C vssd1 vssd1 vccd1 vccd1 _10776_/X sky130_fd_sc_hd__and3_1
X_13564_ _13595_/A _13564_/B _13564_/C vssd1 vssd1 vccd1 vccd1 _13565_/A sky130_fd_sc_hd__and3_1
XFILLER_13_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15303_ _15322_/CLK _15303_/D vssd1 vssd1 vccd1 vccd1 _15303_/Q sky130_fd_sc_hd__dfxtp_1
X_12515_ _15851_/Q _12744_/B _12519_/C vssd1 vssd1 vccd1 vccd1 _12515_/Y sky130_fd_sc_hd__nand3_1
X_16283_ _16283_/CLK _16283_/D vssd1 vssd1 vccd1 vccd1 _16283_/Q sky130_fd_sc_hd__dfxtp_1
X_13495_ _13538_/A _13495_/B _13495_/C vssd1 vssd1 vccd1 vccd1 _13496_/A sky130_fd_sc_hd__and3_1
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15234_ _15259_/CLK _15234_/D vssd1 vssd1 vccd1 vccd1 _15234_/Q sky130_fd_sc_hd__dfxtp_1
X_12446_ _12454_/A _12446_/B _12446_/C vssd1 vssd1 vccd1 vccd1 _12447_/A sky130_fd_sc_hd__and3_1
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ _12377_/A vssd1 vssd1 vccd1 vccd1 _12377_/X sky130_fd_sc_hd__clkbuf_4
X_15165_ _16365_/Q _15165_/B _15165_/C vssd1 vssd1 vccd1 vccd1 _15168_/B sky130_fd_sc_hd__nand3_1
X_11328_ _11326_/B _11326_/C _11327_/X vssd1 vssd1 vccd1 vccd1 _11329_/C sky130_fd_sc_hd__o21ai_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ _16129_/Q _14137_/C _14069_/X vssd1 vssd1 vccd1 vccd1 _14118_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ _16347_/Q _15131_/B _15096_/C vssd1 vssd1 vccd1 vccd1 _15099_/B sky130_fd_sc_hd__nand3_1
XFILLER_141_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11259_ _15655_/Q _11431_/B _11259_/C vssd1 vssd1 vccd1 vccd1 _11268_/B sky130_fd_sc_hd__and3_1
X_14047_ _16115_/Q _14046_/C _14004_/X vssd1 vssd1 vccd1 vccd1 _14048_/B sky130_fd_sc_hd__a21o_1
XFILLER_140_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15998_ _16052_/CLK _15998_/D vssd1 vssd1 vccd1 vccd1 _15998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ _16312_/Q _14953_/C _14789_/X vssd1 vssd1 vccd1 vccd1 _14949_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15337_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08470_ _15314_/Q _15313_/Q _15312_/Q _07608_/X vssd1 vssd1 vccd1 vccd1 _15223_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_23_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09022_ _09022_/A vssd1 vssd1 vccd1 vccd1 _15305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09924_ _09924_/A vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _15435_/Q _09911_/B _09855_/C vssd1 vssd1 vccd1 vccd1 _09855_/Y sky130_fd_sc_hd__nand3_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _08821_/A _08806_/B _08806_/C vssd1 vssd1 vccd1 vccd1 _08807_/A sky130_fd_sc_hd__and3_1
XFILLER_85_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09786_ _10940_/A vssd1 vssd1 vccd1 vccd1 _09786_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08737_ _15263_/Q _08794_/B _08745_/C vssd1 vssd1 vccd1 vccd1 _08742_/A sky130_fd_sc_hd__and3_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15254_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _08667_/B _08667_/C _08541_/X vssd1 vssd1 vccd1 vccd1 _08669_/C sky130_fd_sc_hd__o21ai_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _14071_/B vssd1 vssd1 vccd1 vccd1 _15021_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08599_ _11037_/A vssd1 vssd1 vccd1 vccd1 _08839_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10628_/A _10628_/B _10629_/X vssd1 vssd1 vccd1 vccd1 _15555_/D sky130_fd_sc_hd__a21oi_1
X_10561_ _15546_/Q _10734_/B _10561_/C vssd1 vssd1 vccd1 vccd1 _10572_/A sky130_fd_sc_hd__and3_1
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ _12299_/B _12299_/C _12188_/X vssd1 vssd1 vccd1 vccd1 _12301_/C sky130_fd_sc_hd__o21ai_1
X_13280_ _13272_/B _13273_/C _13276_/X _13278_/Y vssd1 vssd1 vccd1 vccd1 _13281_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10492_ _15534_/Q _10492_/B _10492_/C vssd1 vssd1 vccd1 vccd1 _10492_/Y sky130_fd_sc_hd__nand3_1
XFILLER_108_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ _15806_/Q _12458_/B _12235_/C vssd1 vssd1 vccd1 vccd1 _12231_/Y sky130_fd_sc_hd__nand3_1
XFILLER_135_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12162_ _12170_/A _12162_/B _12162_/C vssd1 vssd1 vccd1 vccd1 _12163_/A sky130_fd_sc_hd__and3_1
XFILLER_107_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11113_ _15633_/Q _11289_/B _11113_/C vssd1 vssd1 vccd1 vccd1 _11113_/X sky130_fd_sc_hd__and3_1
XFILLER_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12093_ _12377_/A vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11044_ _11058_/C vssd1 vssd1 vccd1 vccd1 _11066_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15921_ _07603_/A _15921_/D vssd1 vssd1 vccd1 vccd1 _15921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15852_ _15907_/CLK _15852_/D vssd1 vssd1 vccd1 vccd1 _15852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14803_ _14797_/A _14800_/B _14646_/X vssd1 vssd1 vccd1 vccd1 _14811_/C sky130_fd_sc_hd__o21a_1
XFILLER_18_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15783_ _15794_/CLK _15783_/D vssd1 vssd1 vccd1 vccd1 _15783_/Q sky130_fd_sc_hd__dfxtp_2
X_12995_ _12995_/A vssd1 vssd1 vccd1 vccd1 _15928_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_56_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _16317_/CLK sky130_fd_sc_hd__clkbuf_16
X_14734_ _07710_/X _14733_/A _14614_/X vssd1 vssd1 vccd1 vccd1 _14734_/Y sky130_fd_sc_hd__a21oi_1
X_11946_ _15761_/Q _12174_/B _11950_/C vssd1 vssd1 vccd1 vccd1 _11946_/Y sky130_fd_sc_hd__nand3_1
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14665_ _16248_/Q _14743_/B _14665_/C vssd1 vssd1 vccd1 vccd1 _14668_/B sky130_fd_sc_hd__nand3_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12107_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13616_ _13616_/A vssd1 vssd1 vccd1 vccd1 _16033_/D sky130_fd_sc_hd__clkbuf_1
X_10828_ _10822_/B _10823_/C _10825_/X _10826_/Y vssd1 vssd1 vccd1 vccd1 _10829_/C
+ sky130_fd_sc_hd__a211o_1
X_14596_ _14590_/B _14591_/C _14600_/A _14594_/Y vssd1 vssd1 vccd1 vccd1 _14600_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_71_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16335_ _16344_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 _16335_/Q sky130_fd_sc_hd__dfxtp_2
X_13547_ _13547_/A vssd1 vssd1 vccd1 vccd1 _16021_/D sky130_fd_sc_hd__clkbuf_1
X_10759_ _10792_/C vssd1 vssd1 vccd1 vccd1 _10798_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16266_ _16273_/CLK _16266_/D vssd1 vssd1 vccd1 vccd1 _16266_/Q sky130_fd_sc_hd__dfxtp_1
X_13478_ _16012_/Q _13484_/C _13269_/X vssd1 vssd1 vccd1 vccd1 _13480_/C sky130_fd_sc_hd__a21o_1
X_15217_ _16224_/CLK _15217_/D vssd1 vssd1 vccd1 vccd1 state1[2] sky130_fd_sc_hd__dfxtp_2
X_12429_ _15839_/Q _12434_/C _12370_/X vssd1 vssd1 vccd1 vccd1 _12431_/C sky130_fd_sc_hd__a21o_1
X_16197_ _16222_/CLK _16197_/D vssd1 vssd1 vccd1 vccd1 _16197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15148_ _15146_/A _15146_/B _15147_/X vssd1 vssd1 vccd1 vccd1 _16354_/D sky130_fd_sc_hd__a21oi_1
XFILLER_114_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07970_ _13626_/C _07970_/B vssd1 vssd1 vccd1 vccd1 _07970_/X sky130_fd_sc_hd__or2_1
X_15079_ _15074_/A _15077_/B _15043_/X vssd1 vssd1 vccd1 vccd1 _15085_/C sky130_fd_sc_hd__o21a_1
X_09640_ _15401_/Q _09813_/B _09644_/C vssd1 vssd1 vccd1 vccd1 _09640_/Y sky130_fd_sc_hd__nand3_1
XFILLER_95_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09571_ _15392_/Q _09577_/C _09453_/X vssd1 vssd1 vccd1 vccd1 _09571_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_47_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16189_/CLK sky130_fd_sc_hd__clkbuf_16
X_08522_ _15232_/Q _10963_/C _08522_/C vssd1 vssd1 vccd1 vccd1 _08535_/A sky130_fd_sc_hd__and3_1
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08453_ _08453_/A _08453_/B vssd1 vssd1 vccd1 vccd1 _08453_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08384_ _08384_/A _08384_/B _08384_/C vssd1 vssd1 vccd1 vccd1 _08386_/A sky130_fd_sc_hd__or3_1
XFILLER_51_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09005_ _09011_/A _09002_/Y _09004_/Y _08999_/C vssd1 vssd1 vccd1 vccd1 _09007_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09907_ _09922_/A _09907_/B _09907_/C vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__and3_1
XFILLER_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _15433_/Q _09950_/B _09847_/C vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__and3_1
X_09769_ _15422_/Q vssd1 vssd1 vccd1 vccd1 _09784_/C sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_38_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16114_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11800_ _11801_/B _11801_/C _11801_/A vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__a21o_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12778_/X _12779_/Y _12774_/B _12775_/C vssd1 vssd1 vccd1 vccd1 _12782_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _15736_/Q _15735_/Q _15734_/Q _11560_/X vssd1 vssd1 vccd1 vccd1 _15728_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14446_/Y _14449_/X _14415_/X vssd1 vssd1 vccd1 vccd1 _14450_/Y sky130_fd_sc_hd__a21oi_1
X_11662_ _15718_/Q _11719_/B _11662_/C vssd1 vssd1 vccd1 vccd1 _11670_/B sky130_fd_sc_hd__and3_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _15998_/Q _13605_/B _13401_/C vssd1 vssd1 vccd1 vccd1 _13408_/B sky130_fd_sc_hd__and3_1
X_10613_ _10609_/X _10611_/Y _10612_/Y _10607_/C vssd1 vssd1 vccd1 vccd1 _10615_/B
+ sky130_fd_sc_hd__o211ai_1
X_14381_ _14427_/A _14381_/B _14386_/A vssd1 vssd1 vccd1 vccd1 _16180_/D sky130_fd_sc_hd__nor3_1
X_11593_ _15707_/Q _11599_/C _11472_/X vssd1 vssd1 vccd1 vccd1 _11593_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16120_ _16123_/CLK _16120_/D vssd1 vssd1 vccd1 vccd1 _16120_/Q sky130_fd_sc_hd__dfxtp_1
X_10544_ _10559_/A _10544_/B _10544_/C vssd1 vssd1 vccd1 vccd1 _10545_/A sky130_fd_sc_hd__and3_1
X_13332_ _13332_/A vssd1 vssd1 vccd1 vccd1 _15984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16051_ _16060_/CLK _16051_/D vssd1 vssd1 vccd1 vccd1 _16051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10475_ _15532_/Q _10512_/C _10474_/X vssd1 vssd1 vccd1 vccd1 _10477_/B sky130_fd_sc_hd__a21oi_1
X_13263_ _13276_/C vssd1 vssd1 vccd1 vccd1 _13291_/C sky130_fd_sc_hd__clkbuf_1
X_15002_ _14996_/A _14999_/B _14845_/X vssd1 vssd1 vccd1 vccd1 _15010_/C sky130_fd_sc_hd__o21a_1
X_12214_ _15805_/Q _12383_/B _12216_/C vssd1 vssd1 vccd1 vccd1 _12214_/X sky130_fd_sc_hd__and3_1
X_13194_ _14099_/B vssd1 vssd1 vccd1 vccd1 _13194_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12145_ _15794_/Q _12150_/C _12086_/X vssd1 vssd1 vccd1 vccd1 _12147_/C sky130_fd_sc_hd__a21o_1
XFILLER_123_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12076_ _15788_/Q _15790_/Q _15789_/Q _11847_/X vssd1 vssd1 vccd1 vccd1 _15782_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11027_ _15619_/Q _11143_/B _11027_/C vssd1 vssd1 vccd1 vccd1 _11036_/B sky130_fd_sc_hd__and3_1
X_15904_ _15907_/CLK _15904_/D vssd1 vssd1 vccd1 vccd1 _15904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15835_ _15907_/CLK _15835_/D vssd1 vssd1 vccd1 vccd1 _15835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15766_ _15794_/CLK _15766_/D vssd1 vssd1 vccd1 vccd1 _15766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12978_ _12977_/B _12977_/C _12758_/X vssd1 vssd1 vccd1 vccd1 _12979_/C sky130_fd_sc_hd__o21ai_1
XFILLER_33_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14717_ _16259_/Q _14755_/B _14717_/C vssd1 vssd1 vccd1 vccd1 _14720_/A sky130_fd_sc_hd__and3_1
X_11929_ _15760_/Q _12099_/B _11931_/C vssd1 vssd1 vccd1 vccd1 _11929_/X sky130_fd_sc_hd__and3_1
X_15697_ _15794_/CLK _15697_/D vssd1 vssd1 vccd1 vccd1 _15697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14648_ _14648_/A _14654_/C vssd1 vssd1 vccd1 vccd1 _14648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_17 _14593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _10341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 _13693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14579_ _14579_/A _14579_/B vssd1 vssd1 vccd1 vccd1 _16223_/D sky130_fd_sc_hd__nor2_1
X_16318_ _16327_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 _16318_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16249_ _16268_/CLK _16249_/D vssd1 vssd1 vccd1 vccd1 _16249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07953_ _13523_/C _07918_/B _07952_/X vssd1 vssd1 vccd1 vccd1 _07983_/A sky130_fd_sc_hd__o21ai_4
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07884_ _15620_/Q _07885_/B vssd1 vssd1 vccd1 vccd1 _07886_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09623_ _15399_/Q _09623_/B _09623_/C vssd1 vssd1 vccd1 vccd1 _09623_/Y sky130_fd_sc_hd__nand3_1
X_09554_ _09575_/A _09554_/B _09554_/C vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__and3_1
X_08505_ _15229_/Q _08753_/B _08505_/C vssd1 vssd1 vccd1 vccd1 _08505_/Y sky130_fd_sc_hd__nand3_1
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09485_ _15379_/Q _09528_/C _09316_/X vssd1 vssd1 vccd1 vccd1 _09487_/B sky130_fd_sc_hd__a21oi_1
XFILLER_102_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08436_ _08436_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08436_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08367_ _08272_/A _08272_/B _08329_/A _08366_/X vssd1 vssd1 vccd1 vccd1 _08368_/B
+ sky130_fd_sc_hd__a31o_1
X_08298_ _08298_/A _08341_/A vssd1 vssd1 vccd1 vccd1 _08321_/A sky130_fd_sc_hd__xnor2_2
XFILLER_125_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _10260_/A vssd1 vssd1 vccd1 vccd1 _15498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10191_ _15489_/Q _10363_/B _10191_/C vssd1 vssd1 vccd1 vccd1 _10191_/X sky130_fd_sc_hd__and3_1
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13950_ _16096_/Q _13950_/B _13957_/C vssd1 vssd1 vccd1 vccd1 _13953_/A sky130_fd_sc_hd__and3_1
XFILLER_86_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12901_ _15914_/Q _12954_/B _12908_/C vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__and3_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13881_ _13881_/A _13881_/B _13881_/C vssd1 vssd1 vccd1 vccd1 _13882_/C sky130_fd_sc_hd__nand3_1
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15620_ _15620_/CLK _15620_/D vssd1 vssd1 vccd1 vccd1 _15620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _15903_/Q _12996_/B _12832_/C vssd1 vssd1 vccd1 vccd1 _12832_/X sky130_fd_sc_hd__and3_1
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15655_/CLK _15551_/D vssd1 vssd1 vccd1 vccd1 _15551_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12763_/A vssd1 vssd1 vccd1 vccd1 _12778_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14513_/C vssd1 vssd1 vccd1 vccd1 _14525_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11714_ _15726_/Q _11719_/C _11713_/X vssd1 vssd1 vccd1 vccd1 _11714_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _15483_/CLK _15482_/D vssd1 vssd1 vccd1 vccd1 _15482_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12919_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14433_/A vssd1 vssd1 vccd1 vccd1 _16190_/D sky130_fd_sc_hd__clkbuf_1
X_11645_ _11643_/Y _11639_/C _11641_/X _11642_/Y vssd1 vssd1 vccd1 vccd1 _11646_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14364_ _14364_/A vssd1 vssd1 vccd1 vccd1 _14532_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11576_ _15705_/Q _11576_/B _11576_/C vssd1 vssd1 vccd1 vccd1 _11576_/X sky130_fd_sc_hd__and3_1
XFILLER_11_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16103_ _16103_/CLK _16103_/D vssd1 vssd1 vccd1 vccd1 _16103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13315_ _13341_/C vssd1 vssd1 vccd1 vccd1 _13349_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10527_ _10527_/A vssd1 vssd1 vccd1 vccd1 _10540_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14295_ _14295_/A _14295_/B _14295_/C vssd1 vssd1 vccd1 vccd1 _14296_/C sky130_fd_sc_hd__nand3_1
XFILLER_109_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16034_ _16052_/CLK _16034_/D vssd1 vssd1 vccd1 vccd1 _16034_/Q sky130_fd_sc_hd__dfxtp_1
X_10458_ _10629_/A _10463_/C vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__or2_1
XFILLER_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13246_ _15971_/Q _13349_/B _13246_/C vssd1 vssd1 vccd1 vccd1 _13255_/B sky130_fd_sc_hd__and3_1
X_10389_ _15519_/Q _10446_/B _10389_/C vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__and3_1
X_13177_ _13177_/A vssd1 vssd1 vccd1 vccd1 _15957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12128_ _12126_/A _12126_/B _12127_/X vssd1 vssd1 vccd1 vccd1 _15789_/D sky130_fd_sc_hd__a21oi_1
X_12059_ _12057_/Y _12053_/C _12066_/A _12056_/Y vssd1 vssd1 vccd1 vccd1 _12066_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15818_ _15818_/CLK _15818_/D vssd1 vssd1 vccd1 vccd1 _15818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15749_ _15794_/CLK _15749_/D vssd1 vssd1 vccd1 vccd1 _15749_/Q sky130_fd_sc_hd__dfxtp_1
X_09270_ _15346_/Q _09496_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09270_/X sky130_fd_sc_hd__and3_1
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08221_ _08221_/A _08289_/A vssd1 vssd1 vccd1 vccd1 _08259_/A sky130_fd_sc_hd__xnor2_4
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08152_ _15306_/Q _08152_/B vssd1 vssd1 vccd1 vccd1 _08152_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08083_ _08083_/A _07781_/B vssd1 vssd1 vccd1 vccd1 _08083_/X sky130_fd_sc_hd__or2b_1
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _08999_/A _08985_/B _08985_/C vssd1 vssd1 vccd1 vccd1 _08986_/A sky130_fd_sc_hd__and3_1
XFILLER_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07936_ _15270_/Q _08156_/B vssd1 vssd1 vccd1 vccd1 _07937_/B sky130_fd_sc_hd__xnor2_1
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07867_ _14117_/C _08012_/B vssd1 vssd1 vccd1 vccd1 _07868_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _15397_/Q _09644_/C _09605_/X vssd1 vssd1 vccd1 vccd1 _09608_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07798_ _12874_/A _08077_/B vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__xnor2_1
XFILLER_73_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09537_ _09708_/A _09537_/B _09537_/C vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__or3_1
X_09468_ _15376_/Q _09466_/C _09467_/X vssd1 vssd1 vccd1 vccd1 _09469_/B sky130_fd_sc_hd__a21oi_1
X_08419_ _08420_/A spike_out[0] _08420_/C vssd1 vssd1 vccd1 vccd1 _08421_/B sky130_fd_sc_hd__o21a_1
X_09399_ _09396_/X _09397_/Y _09398_/Y _09394_/C vssd1 vssd1 vccd1 vccd1 _09401_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ _11509_/A _11430_/B _11434_/B vssd1 vssd1 vccd1 vccd1 _15680_/D sky130_fd_sc_hd__nor3_1
XFILLER_11_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _15671_/Q _11367_/C _11184_/X vssd1 vssd1 vccd1 vccd1 _11361_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10312_ _15507_/Q _10492_/B _10312_/C vssd1 vssd1 vccd1 vccd1 _10312_/Y sky130_fd_sc_hd__nand3_1
X_13100_ _13679_/A vssd1 vssd1 vccd1 vccd1 _14291_/A sky130_fd_sc_hd__buf_2
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11292_ _11286_/B _11287_/C _11289_/X _11290_/Y vssd1 vssd1 vccd1 vccd1 _11293_/C
+ sky130_fd_sc_hd__a211o_1
X_14080_ _16121_/Q _14080_/B _14080_/C vssd1 vssd1 vccd1 vccd1 _14080_/X sky130_fd_sc_hd__and3_1
X_10243_ _10244_/B _10244_/C _10244_/A vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__a21o_1
X_13031_ _13151_/A _13031_/B _13031_/C vssd1 vssd1 vccd1 vccd1 _13033_/B sky130_fd_sc_hd__or3_1
XFILLER_98_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10174_ _10210_/A _10174_/B _10174_/C vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__and3_1
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14982_ _16320_/Q _14981_/C _14942_/X vssd1 vssd1 vccd1 vccd1 _14984_/C sky130_fd_sc_hd__a21o_1
X_13933_ _16106_/Q _16105_/Q _16104_/Q _13723_/X vssd1 vssd1 vccd1 vccd1 _16089_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13864_ _13864_/A vssd1 vssd1 vccd1 vccd1 _16078_/D sky130_fd_sc_hd__clkbuf_1
X_15603_ _15194_/Q _15603_/D vssd1 vssd1 vccd1 vccd1 _15603_/Q sky130_fd_sc_hd__dfxtp_2
X_12815_ _12851_/A _12815_/B _12815_/C vssd1 vssd1 vccd1 vccd1 _12816_/A sky130_fd_sc_hd__and3_1
X_13795_ _13792_/X _13793_/Y _13794_/Y _13789_/C vssd1 vssd1 vccd1 vccd1 _13797_/B
+ sky130_fd_sc_hd__o211ai_1
X_15534_ _15655_/CLK _15534_/D vssd1 vssd1 vccd1 vccd1 _15534_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _12744_/Y _12740_/C _12751_/A _12743_/Y vssd1 vssd1 vccd1 vccd1 _12751_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ _15484_/CLK _15465_/D vssd1 vssd1 vccd1 vccd1 _15465_/Q sky130_fd_sc_hd__dfxtp_1
X_12677_ _15877_/Q _12793_/B _12684_/C vssd1 vssd1 vccd1 vccd1 _12677_/Y sky130_fd_sc_hd__nand3_1
XFILLER_129_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14416_ _14368_/X _14411_/B _14415_/X vssd1 vssd1 vccd1 vccd1 _14416_/Y sky130_fd_sc_hd__a21oi_1
X_11628_ _15713_/Q _11797_/B _11635_/C vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__nand3_1
X_15396_ _15483_/CLK _15396_/D vssd1 vssd1 vccd1 vccd1 _15396_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14347_ _14352_/A _14346_/Y _14342_/B _14343_/C vssd1 vssd1 vccd1 vccd1 _14349_/B
+ sky130_fd_sc_hd__o211a_1
X_11559_ _11559_/A vssd1 vssd1 vccd1 vccd1 _15700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ _14190_/X _14276_/B _14277_/Y vssd1 vssd1 vccd1 vccd1 _16158_/D sky130_fd_sc_hd__o21a_1
X_16017_ _16040_/CLK _16017_/D vssd1 vssd1 vccd1 vccd1 _16017_/Q sky130_fd_sc_hd__dfxtp_2
X_13229_ _13222_/B _13223_/C _13226_/X _13227_/Y vssd1 vssd1 vccd1 vccd1 _13230_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08770_ _15268_/Q _08775_/C _08524_/X vssd1 vssd1 vccd1 vccd1 _08770_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07721_ _15225_/Q _15223_/Q vssd1 vssd1 vccd1 vccd1 _08125_/B sky130_fd_sc_hd__xor2_2
XFILLER_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07652_ _07638_/B _07639_/C _07666_/A _07650_/Y vssd1 vssd1 vccd1 vccd1 _07666_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_19_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09322_ _09323_/B _09323_/C _09323_/A vssd1 vssd1 vccd1 vccd1 _09324_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09253_ _09288_/A _09253_/B _09253_/C vssd1 vssd1 vccd1 vccd1 _09254_/A sky130_fd_sc_hd__and3_1
X_08204_ _08081_/A _08081_/B _08203_/X vssd1 vssd1 vccd1 vccd1 _08220_/A sky130_fd_sc_hd__a21bo_1
X_09184_ _09184_/A _09184_/B vssd1 vssd1 vccd1 vccd1 _09190_/C sky130_fd_sc_hd__nor2_1
XFILLER_119_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08135_ _08241_/A _08241_/B vssd1 vssd1 vccd1 vccd1 _08252_/A sky130_fd_sc_hd__xnor2_4
XFILLER_147_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08066_ _14627_/C _08066_/B vssd1 vssd1 vccd1 vccd1 _08066_/X sky130_fd_sc_hd__or2_1
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08968_ _08989_/C vssd1 vssd1 vccd1 vccd1 _09001_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07919_ _13420_/C _07952_/B vssd1 vssd1 vccd1 vccd1 _07920_/B sky130_fd_sc_hd__xnor2_4
X_08899_ _08942_/A _08899_/B _08899_/C vssd1 vssd1 vccd1 vccd1 _08900_/A sky130_fd_sc_hd__and3_1
XFILLER_72_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930_ _15604_/Q _10939_/B _13474_/A vssd1 vssd1 vccd1 vccd1 _10936_/A sky130_fd_sc_hd__and3_1
XFILLER_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861_ _10859_/A _10859_/B _10860_/X vssd1 vssd1 vccd1 vccd1 _15591_/D sky130_fd_sc_hd__a21oi_1
XFILLER_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12600_/A vssd1 vssd1 vccd1 vccd1 _15865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13580_/A _13580_/B _13580_/C vssd1 vssd1 vccd1 vccd1 _13581_/C sky130_fd_sc_hd__nand3_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _15582_/Q _11078_/B _10792_/C vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__and3_1
XFILLER_52_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _15862_/Q _15861_/Q _15860_/Q _12418_/X vssd1 vssd1 vccd1 vccd1 _15854_/D
+ sky130_fd_sc_hd__o31a_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _15259_/CLK _15250_/D vssd1 vssd1 vccd1 vccd1 _15250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12462_ _15844_/Q _12575_/B _12462_/C vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__and3_1
XFILLER_149_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14201_ _14201_/A _14201_/B vssd1 vssd1 vccd1 vccd1 _16142_/D sky130_fd_sc_hd__nor2_1
XFILLER_138_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11413_ _11413_/A vssd1 vssd1 vccd1 vccd1 _15678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15181_ _15181_/A _15181_/B vssd1 vssd1 vccd1 vccd1 _15181_/X sky130_fd_sc_hd__or2_1
X_12393_ _15832_/Q _12507_/B _12399_/C vssd1 vssd1 vccd1 vccd1 _12393_/Y sky130_fd_sc_hd__nand3_1
XFILLER_138_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _14132_/A _14132_/B vssd1 vssd1 vccd1 vccd1 _14132_/Y sky130_fd_sc_hd__nor2_1
X_11344_ _11365_/A _11344_/B _11344_/C vssd1 vssd1 vccd1 vccd1 _11345_/A sky130_fd_sc_hd__and3_1
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14063_ _14063_/A _14063_/B vssd1 vssd1 vccd1 vccd1 _16115_/D sky130_fd_sc_hd__nor2_1
XFILLER_125_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11275_/A vssd1 vssd1 vccd1 vccd1 _11289_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13014_ _13014_/A _13014_/B _13014_/C vssd1 vssd1 vccd1 vccd1 _13015_/A sky130_fd_sc_hd__and3_1
X_10226_ _10224_/A _10224_/B _10225_/X vssd1 vssd1 vccd1 vccd1 _15492_/D sky130_fd_sc_hd__a21oi_1
XFILLER_67_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10157_ _10736_/A vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_121_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ _10097_/A _10088_/B _10088_/C vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__and3_1
XFILLER_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14965_ _14964_/X _14967_/C _14893_/X vssd1 vssd1 vccd1 vccd1 _14966_/B sky130_fd_sc_hd__o21ai_1
XFILLER_48_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13916_ _15186_/A _13916_/B vssd1 vssd1 vccd1 vccd1 _13917_/B sky130_fd_sc_hd__and2_1
XFILLER_62_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14896_ _14772_/X _14895_/A _14815_/X vssd1 vssd1 vccd1 vccd1 _14896_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _13847_/A vssd1 vssd1 vccd1 vccd1 _14270_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13778_ _13852_/A _13778_/B _13782_/A vssd1 vssd1 vccd1 vccd1 _16063_/D sky130_fd_sc_hd__nor3_1
X_15517_ _15655_/CLK _15517_/D vssd1 vssd1 vccd1 vccd1 _15517_/Q sky130_fd_sc_hd__dfxtp_1
X_12729_ _15885_/Q _12840_/B _12729_/C vssd1 vssd1 vccd1 vccd1 _12729_/Y sky130_fd_sc_hd__nand3_1
XFILLER_148_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15448_ _15484_/CLK _15448_/D vssd1 vssd1 vccd1 vccd1 _15448_/Q sky130_fd_sc_hd__dfxtp_1
X_15379_ _15484_/CLK _15379_/D vssd1 vssd1 vccd1 vccd1 _15379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09940_ _09939_/B _09939_/C _09884_/X vssd1 vssd1 vccd1 vccd1 _09941_/C sky130_fd_sc_hd__o21ai_1
X_09871_ _09877_/A _09868_/Y _09870_/Y _09865_/C vssd1 vssd1 vccd1 vccd1 _09873_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08822_ _08822_/A vssd1 vssd1 vccd1 vccd1 _15275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08753_ _15265_/Q _08753_/B _08753_/C vssd1 vssd1 vccd1 vccd1 _08753_/Y sky130_fd_sc_hd__nand3_1
XFILLER_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ input8/X vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__buf_4
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08684_ _08684_/A vssd1 vssd1 vccd1 vccd1 _15254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ _14980_/A vssd1 vssd1 vccd1 vccd1 _15165_/B sky130_fd_sc_hd__clkbuf_4
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09305_ _09536_/A vssd1 vssd1 vccd1 vccd1 _09345_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09236_ _15340_/Q _09290_/B _09236_/C vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__and3_1
X_09167_ _15330_/Q _09173_/C _09166_/X vssd1 vssd1 vccd1 vccd1 _09167_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08118_ _15333_/Q vssd1 vssd1 vccd1 vccd1 _09256_/A sky130_fd_sc_hd__inv_2
XFILLER_119_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _09096_/X _09097_/Y _09093_/B _09094_/C vssd1 vssd1 vccd1 vccd1 _09100_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_134_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08049_ _15845_/Q _08049_/B vssd1 vssd1 vccd1 vccd1 _08049_/Y sky130_fd_sc_hd__nand2_1
X_11060_ _11058_/X _11059_/Y _11054_/B _11055_/C vssd1 vssd1 vccd1 vccd1 _11062_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_89_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10011_ _15461_/Q _10016_/C _09778_/X vssd1 vssd1 vccd1 vccd1 _10013_/C sky130_fd_sc_hd__a21o_1
XFILLER_135_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14750_ _16267_/Q _14833_/B _14755_/C vssd1 vssd1 vccd1 vccd1 _14758_/A sky130_fd_sc_hd__and3_1
X_11962_ _15772_/Q _15771_/Q _15770_/Q _11847_/X vssd1 vssd1 vccd1 vccd1 _15764_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_57_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13701_ _16051_/Q _14093_/B _13701_/C vssd1 vssd1 vccd1 vccd1 _13711_/A sky130_fd_sc_hd__and3_1
X_10913_ _10920_/B _10913_/B vssd1 vssd1 vccd1 vccd1 _10915_/A sky130_fd_sc_hd__or2_1
X_14681_ _14879_/A vssd1 vssd1 vccd1 vccd1 _14843_/A sky130_fd_sc_hd__clkbuf_2
X_11893_ _11901_/B _11893_/B vssd1 vssd1 vccd1 vccd1 _11895_/A sky130_fd_sc_hd__or2_1
X_13632_ _13664_/A _13632_/B _13632_/C vssd1 vssd1 vccd1 vccd1 _13633_/A sky130_fd_sc_hd__and3_1
XFILLER_72_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ _10842_/Y _10838_/C _10840_/X _10841_/Y vssd1 vssd1 vccd1 vccd1 _10845_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16377__26 vssd1 vssd1 vccd1 vccd1 _16377__26/HI io_oeb[9] sky130_fd_sc_hd__conb_1
X_16351_ _16358_/CLK _16351_/D vssd1 vssd1 vccd1 vccd1 _16351_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13563_ _13561_/B _13561_/C _13562_/X vssd1 vssd1 vccd1 vccd1 _13564_/C sky130_fd_sc_hd__o21ai_1
X_10775_ _10775_/A vssd1 vssd1 vccd1 vccd1 _15578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15302_ _15322_/CLK _15302_/D vssd1 vssd1 vccd1 vccd1 _15302_/Q sky130_fd_sc_hd__dfxtp_1
X_12514_ _13847_/A vssd1 vssd1 vccd1 vccd1 _12744_/B sky130_fd_sc_hd__buf_2
X_16282_ _16283_/CLK _16282_/D vssd1 vssd1 vccd1 vccd1 _16282_/Q sky130_fd_sc_hd__dfxtp_2
X_13494_ _13492_/Y _13488_/C _13490_/X _13491_/Y vssd1 vssd1 vccd1 vccd1 _13495_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15233_ _15254_/CLK _15233_/D vssd1 vssd1 vccd1 vccd1 _15233_/Q sky130_fd_sc_hd__dfxtp_1
X_12445_ _12443_/Y _12438_/C _12441_/X _12442_/Y vssd1 vssd1 vccd1 vccd1 _12446_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15164_ _15175_/A _15164_/B _15168_/A vssd1 vssd1 vccd1 vccd1 _16360_/D sky130_fd_sc_hd__nor3_1
X_12376_ _15831_/Q _12434_/B _12376_/C vssd1 vssd1 vccd1 vccd1 _12376_/X sky130_fd_sc_hd__and3_1
X_14115_ _14125_/C vssd1 vssd1 vccd1 vccd1 _14137_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11327_ _12188_/A vssd1 vssd1 vccd1 vccd1 _11327_/X sky130_fd_sc_hd__clkbuf_2
X_15095_ _15106_/A _15095_/B _15099_/A vssd1 vssd1 vccd1 vccd1 _16342_/D sky130_fd_sc_hd__nor3_1
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14046_ _16115_/Q _14137_/B _14046_/C vssd1 vssd1 vccd1 vccd1 _14046_/X sky130_fd_sc_hd__and3_1
X_11258_ _11373_/A _11258_/B _11262_/B vssd1 vssd1 vccd1 vccd1 _15653_/D sky130_fd_sc_hd__nor3_1
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10209_ _10207_/Y _10202_/C _10204_/X _10205_/Y vssd1 vssd1 vccd1 vccd1 _10210_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_67_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11189_ _11189_/A _11189_/B _11189_/C vssd1 vssd1 vccd1 vccd1 _11190_/A sky130_fd_sc_hd__and3_1
XFILLER_94_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15997_ _16052_/CLK _15997_/D vssd1 vssd1 vccd1 vccd1 _15997_/Q sky130_fd_sc_hd__dfxtp_1
X_14948_ _16312_/Q _15031_/B _14953_/C vssd1 vssd1 vccd1 vccd1 _14956_/A sky130_fd_sc_hd__and3_1
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14879_ _14879_/A vssd1 vssd1 vccd1 vccd1 _15041_/A sky130_fd_sc_hd__buf_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09021_ _09058_/A _09021_/B _09021_/C vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__and3_1
XFILLER_117_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09923_ _09923_/A vssd1 vssd1 vccd1 vccd1 _15445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09854_ _15436_/Q _09855_/C _09794_/X vssd1 vssd1 vccd1 vccd1 _09854_/Y sky130_fd_sc_hd__a21oi_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _08799_/B _08800_/C _08802_/X _08803_/Y vssd1 vssd1 vccd1 vccd1 _08806_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _11229_/A vssd1 vssd1 vccd1 vccd1 _10940_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08736_ _15263_/Q _08775_/C _08735_/X vssd1 vssd1 vccd1 vccd1 _08738_/B sky130_fd_sc_hd__a21oi_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _08839_/A _08667_/B _08667_/C vssd1 vssd1 vccd1 vccd1 _08669_/B sky130_fd_sc_hd__or3_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _13043_/B vssd1 vssd1 vccd1 vccd1 _14071_/B sky130_fd_sc_hd__buf_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ input8/X vssd1 vssd1 vccd1 vccd1 _11037_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ _10560_/A vssd1 vssd1 vccd1 vccd1 _15544_/D sky130_fd_sc_hd__clkbuf_1
X_09219_ _15338_/Q _09444_/B _09222_/C vssd1 vssd1 vccd1 vccd1 _09219_/X sky130_fd_sc_hd__and3_1
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10491_ _15535_/Q _10492_/C _10373_/X vssd1 vssd1 vccd1 vccd1 _10491_/Y sky130_fd_sc_hd__a21oi_1
X_12230_ _12230_/A vssd1 vssd1 vccd1 vccd1 _12458_/B sky130_fd_sc_hd__buf_2
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ _12159_/Y _12154_/C _12157_/X _12158_/Y vssd1 vssd1 vccd1 vccd1 _12162_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _11112_/A vssd1 vssd1 vccd1 vccd1 _15631_/D sky130_fd_sc_hd__clkbuf_1
X_12092_ _15786_/Q _12150_/B _12092_/C vssd1 vssd1 vccd1 vccd1 _12092_/X sky130_fd_sc_hd__and3_1
XFILLER_104_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11043_ _15620_/Q vssd1 vssd1 vccd1 vccd1 _11058_/C sky130_fd_sc_hd__inv_2
X_15920_ _07603_/A _15920_/D vssd1 vssd1 vccd1 vccd1 _15920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15851_ _15907_/CLK _15851_/D vssd1 vssd1 vccd1 vccd1 _15851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14802_ _15001_/A vssd1 vssd1 vccd1 vccd1 _14802_/X sky130_fd_sc_hd__buf_2
X_15782_ _15890_/CLK _15782_/D vssd1 vssd1 vccd1 vccd1 _15782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12994_ _13014_/A _12994_/B _12994_/C vssd1 vssd1 vccd1 vccd1 _12995_/A sky130_fd_sc_hd__and3_1
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14733_ _14733_/A _14733_/B vssd1 vssd1 vccd1 vccd1 _16258_/D sky130_fd_sc_hd__nor2_1
XFILLER_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ _12230_/A vssd1 vssd1 vccd1 vccd1 _12174_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14664_ _14716_/A _14664_/B _14668_/A vssd1 vssd1 vccd1 vccd1 _16243_/D sky130_fd_sc_hd__nor3_1
XFILLER_33_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11876_ _11876_/A vssd1 vssd1 vccd1 vccd1 _15750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13615_ _13664_/A _13615_/B _13615_/C vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__and3_1
X_10827_ _10825_/X _10826_/Y _10822_/B _10823_/C vssd1 vssd1 vccd1 vccd1 _10829_/B
+ sky130_fd_sc_hd__o211ai_1
X_14595_ _14600_/A _14594_/Y _14590_/B _14591_/C vssd1 vssd1 vccd1 vccd1 _14597_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16334_ _16344_/CLK _16334_/D vssd1 vssd1 vccd1 vccd1 _16334_/Q sky130_fd_sc_hd__dfxtp_2
X_13546_ _13595_/A _13546_/B _13546_/C vssd1 vssd1 vccd1 vccd1 _13547_/A sky130_fd_sc_hd__and3_1
X_10758_ _10778_/C vssd1 vssd1 vccd1 vccd1 _10792_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16265_ _16268_/CLK _16265_/D vssd1 vssd1 vccd1 vccd1 _16265_/Q sky130_fd_sc_hd__dfxtp_1
X_13477_ _16012_/Q _13628_/B _13484_/C vssd1 vssd1 vccd1 vccd1 _13480_/B sky130_fd_sc_hd__nand3_1
X_10689_ _11551_/A vssd1 vssd1 vccd1 vccd1 _10916_/A sky130_fd_sc_hd__buf_2
X_15216_ _16367_/CLK _15216_/D vssd1 vssd1 vccd1 vccd1 state1[1] sky130_fd_sc_hd__dfxtp_2
XFILLER_145_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12428_ _15839_/Q _12653_/B _12434_/C vssd1 vssd1 vccd1 vccd1 _12431_/B sky130_fd_sc_hd__nand3_1
X_16196_ _16204_/CLK _16196_/D vssd1 vssd1 vccd1 vccd1 _16196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ _15181_/A _15147_/B vssd1 vssd1 vccd1 vccd1 _15147_/X sky130_fd_sc_hd__or2_1
XFILLER_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12359_ _12359_/A vssd1 vssd1 vccd1 vccd1 _15826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15078_ _15076_/A _15076_/B _15077_/X vssd1 vssd1 vccd1 vccd1 _16336_/D sky130_fd_sc_hd__a21oi_1
XFILLER_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14029_ _14029_/A _14029_/B _14029_/C vssd1 vssd1 vccd1 vccd1 _14030_/A sky130_fd_sc_hd__and3_1
XFILLER_67_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09570_ _15392_/Q _09740_/B _09577_/C vssd1 vssd1 vccd1 vccd1 _09570_/X sky130_fd_sc_hd__and3_1
XFILLER_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08521_ _11424_/A vssd1 vssd1 vccd1 vccd1 _10963_/C sky130_fd_sc_hd__buf_2
XFILLER_24_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08452_ _08462_/B _08452_/B vssd1 vssd1 vccd1 vccd1 _08453_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08383_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08386_/C sky130_fd_sc_hd__nand2_1
XFILLER_149_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09004_ _15303_/Q _09238_/B _09008_/C vssd1 vssd1 vccd1 vccd1 _09004_/Y sky130_fd_sc_hd__nand3_1
XFILLER_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09906_ _09900_/B _09901_/C _09903_/X _09904_/Y vssd1 vssd1 vccd1 vccd1 _09907_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _15433_/Q _09874_/C _09605_/X vssd1 vssd1 vccd1 vccd1 _09839_/B sky130_fd_sc_hd__a21oi_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09768_ _15430_/Q _15429_/Q _15428_/Q _09541_/X vssd1 vssd1 vccd1 vccd1 _15422_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_100_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08719_/A _08719_/B vssd1 vssd1 vccd1 vccd1 _08724_/C sky130_fd_sc_hd__nor2_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09699_/A vssd1 vssd1 vccd1 vccd1 _09931_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _11730_/A vssd1 vssd1 vccd1 vccd1 _15727_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11661_/A _11661_/B _11665_/B vssd1 vssd1 vccd1 vccd1 _15716_/D sky130_fd_sc_hd__nor3_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _13654_/A vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__clkbuf_2
X_10612_ _15553_/Q _10729_/B _10617_/C vssd1 vssd1 vccd1 vccd1 _10612_/Y sky130_fd_sc_hd__nand3_1
X_14380_ _16183_/Q _14546_/B _14380_/C vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__and3_1
X_11592_ _15707_/Q _11819_/B _11599_/C vssd1 vssd1 vccd1 vccd1 _11592_/X sky130_fd_sc_hd__and3_1
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _13339_/A _13331_/B _13331_/C vssd1 vssd1 vccd1 vccd1 _13332_/A sky130_fd_sc_hd__and3_1
XFILLER_128_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10543_ _10537_/B _10538_/C _10540_/X _10541_/Y vssd1 vssd1 vccd1 vccd1 _10544_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16050_ _16050_/CLK _16050_/D vssd1 vssd1 vccd1 vccd1 _16050_/Q sky130_fd_sc_hd__dfxtp_1
X_13262_ _13266_/C vssd1 vssd1 vccd1 vccd1 _13276_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10474_ _11624_/A vssd1 vssd1 vccd1 vccd1 _10474_/X sky130_fd_sc_hd__buf_2
X_15001_ _15001_/A vssd1 vssd1 vccd1 vccd1 _15001_/X sky130_fd_sc_hd__buf_2
X_12213_ _12213_/A vssd1 vssd1 vccd1 vccd1 _15803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ _15962_/Q _13349_/B _13193_/C vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__and3_1
XFILLER_135_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12144_ _15794_/Q _12369_/B _12150_/C vssd1 vssd1 vccd1 vccd1 _12147_/B sky130_fd_sc_hd__nand3_1
XFILLER_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12075_ _12075_/A vssd1 vssd1 vccd1 vccd1 _15781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11026_ _11085_/A _11026_/B _11030_/B vssd1 vssd1 vccd1 vccd1 _15617_/D sky130_fd_sc_hd__nor3_1
X_15903_ _15907_/CLK _15903_/D vssd1 vssd1 vccd1 vccd1 _15903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15834_ _15907_/CLK _15834_/D vssd1 vssd1 vccd1 vccd1 _15834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15765_ _15794_/CLK _15765_/D vssd1 vssd1 vccd1 vccd1 _15765_/Q sky130_fd_sc_hd__dfxtp_2
X_12977_ _13151_/A _12977_/B _12977_/C vssd1 vssd1 vccd1 vccd1 _12979_/B sky130_fd_sc_hd__or3_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11928_ _11928_/A vssd1 vssd1 vccd1 vccd1 _15758_/D sky130_fd_sc_hd__clkbuf_1
X_14716_ _14716_/A _14716_/B _14721_/B vssd1 vssd1 vccd1 vccd1 _16254_/D sky130_fd_sc_hd__nor3_1
XFILLER_33_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15696_ _15763_/CLK _15696_/D vssd1 vssd1 vccd1 vccd1 _15696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14647_ _14641_/A _14644_/B _14646_/X vssd1 vssd1 vccd1 vccd1 _14654_/C sky130_fd_sc_hd__o21a_1
XFILLER_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11859_ _11860_/B _11860_/C _11860_/A vssd1 vssd1 vccd1 vccd1 _11861_/B sky130_fd_sc_hd__a21o_1
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_18 hold24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 _12100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ _14368_/A _08541_/X _14573_/B _14459_/X vssd1 vssd1 vccd1 vccd1 _14579_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13529_ _13529_/A _13529_/B _13529_/C vssd1 vssd1 vccd1 vccd1 _13530_/C sky130_fd_sc_hd__nand3_1
X_16317_ _16317_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 _16317_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16248_ _16268_/CLK _16248_/D vssd1 vssd1 vccd1 vccd1 _16248_/Q sky130_fd_sc_hd__dfxtp_1
X_16179_ _16222_/CLK _16179_/D vssd1 vssd1 vccd1 vccd1 _16179_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07952_ _13420_/C _07952_/B vssd1 vssd1 vccd1 vccd1 _07952_/X sky130_fd_sc_hd__or2_1
XFILLER_141_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07883_ _08016_/A _07883_/B vssd1 vssd1 vccd1 vccd1 _07885_/B sky130_fd_sc_hd__xnor2_4
X_09622_ _15400_/Q _09623_/C _09506_/X vssd1 vssd1 vccd1 vccd1 _09622_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09553_ _09553_/A _09553_/B _09553_/C vssd1 vssd1 vccd1 vccd1 _09554_/C sky130_fd_sc_hd__nand3_1
X_08504_ _13534_/A vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__buf_2
X_09484_ _09522_/C vssd1 vssd1 vccd1 vccd1 _09528_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08435_ _08444_/A _08444_/B vssd1 vssd1 vccd1 vccd1 _08435_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_12_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08366_ _08365_/Y _08271_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08366_/X sky130_fd_sc_hd__o21ba_1
X_08297_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08341_/A sky130_fd_sc_hd__xnor2_1
XFILLER_149_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10190_ _10190_/A vssd1 vssd1 vccd1 vccd1 _15487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12900_ _12900_/A vssd1 vssd1 vccd1 vccd1 _15912_/D sky130_fd_sc_hd__clkbuf_1
X_13880_ _13881_/B _13881_/C _13881_/A vssd1 vssd1 vccd1 vccd1 _13882_/B sky130_fd_sc_hd__a21o_1
X_12831_ _12831_/A vssd1 vssd1 vccd1 vccd1 _15901_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15550_ _15655_/CLK _15550_/D vssd1 vssd1 vccd1 vccd1 _15550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _15896_/Q _15898_/Q _15897_/Q _12704_/X vssd1 vssd1 vccd1 vccd1 _15890_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14505_/C vssd1 vssd1 vccd1 vccd1 _14513_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11713_ _12569_/A vssd1 vssd1 vccd1 vccd1 _11713_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15224_/Q _15481_/D vssd1 vssd1 vccd1 vccd1 _15481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _12695_/B sky130_fd_sc_hd__nor2_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14552_/A _14432_/B _14432_/C vssd1 vssd1 vccd1 vccd1 _14433_/A sky130_fd_sc_hd__and3_1
X_11644_ _11641_/X _11642_/Y _11643_/Y _11639_/C vssd1 vssd1 vccd1 vccd1 _11646_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14363_ _14363_/A vssd1 vssd1 vccd1 vccd1 _14533_/A sky130_fd_sc_hd__clkbuf_2
X_11575_ _11575_/A vssd1 vssd1 vccd1 vccd1 _15703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16102_ _16119_/CLK _16102_/D vssd1 vssd1 vccd1 vccd1 _16102_/Q sky130_fd_sc_hd__dfxtp_1
X_13314_ _13327_/C vssd1 vssd1 vccd1 vccd1 _13341_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_128_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10526_ _11099_/A vssd1 vssd1 vccd1 vccd1 _10645_/A sky130_fd_sc_hd__buf_2
X_14294_ _14295_/B _14295_/C _14295_/A vssd1 vssd1 vccd1 vccd1 _14296_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16033_ _16052_/CLK _16033_/D vssd1 vssd1 vccd1 vccd1 _16033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13245_ _13348_/A _13245_/B _13249_/B vssd1 vssd1 vccd1 vccd1 _15968_/D sky130_fd_sc_hd__nor3_1
X_10457_ _10457_/A _10457_/B vssd1 vssd1 vccd1 vccd1 _10463_/C sky130_fd_sc_hd__nor2_1
XFILLER_124_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13176_ _13223_/A _13176_/B _13176_/C vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__and3_1
X_10388_ _10388_/A vssd1 vssd1 vccd1 vccd1 _10511_/A sky130_fd_sc_hd__buf_2
XFILLER_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ _12352_/A _12130_/C vssd1 vssd1 vccd1 vccd1 _12127_/X sky130_fd_sc_hd__or2_1
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12058_ _12066_/A _12056_/Y _12057_/Y _12053_/C vssd1 vssd1 vccd1 vccd1 _12060_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11009_ _11006_/X _11007_/Y _11008_/Y _11003_/C vssd1 vssd1 vccd1 vccd1 _11011_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15817_ _15907_/CLK _15817_/D vssd1 vssd1 vccd1 vccd1 _15817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15748_ _15794_/CLK _15748_/D vssd1 vssd1 vccd1 vccd1 _15748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15679_ _15763_/CLK _15679_/D vssd1 vssd1 vccd1 vccd1 _15679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08220_ _08220_/A _08220_/B vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__xnor2_2
XFILLER_61_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08151_ _08151_/A _08151_/B vssd1 vssd1 vccd1 vccd1 _08175_/A sky130_fd_sc_hd__xnor2_4
X_08082_ _08082_/A _08203_/A vssd1 vssd1 vccd1 vccd1 _08143_/A sky130_fd_sc_hd__xnor2_4
XFILLER_134_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08984_ _08976_/B _08977_/C _08981_/X _08982_/Y vssd1 vssd1 vccd1 vccd1 _08985_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_130_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07935_ _07935_/A _07935_/B vssd1 vssd1 vccd1 vccd1 _08156_/B sky130_fd_sc_hd__xor2_4
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07866_ _15999_/Q _08007_/B vssd1 vssd1 vccd1 vccd1 _08012_/B sky130_fd_sc_hd__xnor2_2
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09605_ _10181_/A vssd1 vssd1 vccd1 vccd1 _09605_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07797_ _14546_/C _07797_/B vssd1 vssd1 vccd1 vccd1 _08077_/B sky130_fd_sc_hd__xnor2_2
X_09536_ _09536_/A vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09467_ _10044_/A vssd1 vssd1 vccd1 vccd1 _09467_/X sky130_fd_sc_hd__buf_2
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08418_ state1[1] vssd1 vssd1 vccd1 vccd1 _08420_/A sky130_fd_sc_hd__inv_2
X_09398_ _15364_/Q _09572_/B _09403_/C vssd1 vssd1 vccd1 vccd1 _09398_/Y sky130_fd_sc_hd__nand3_1
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08349_ _08349_/A _08349_/B _08349_/C vssd1 vssd1 vccd1 vccd1 _08350_/B sky130_fd_sc_hd__nand3_1
XFILLER_137_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _15671_/Q _11533_/B _11367_/C vssd1 vssd1 vccd1 vccd1 _11360_/X sky130_fd_sc_hd__and3_1
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10311_ _15508_/Q _10312_/C _10083_/X vssd1 vssd1 vccd1 vccd1 _10311_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11291_ _11289_/X _11290_/Y _11286_/B _11287_/C vssd1 vssd1 vccd1 vccd1 _11293_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_98_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13030_ _13283_/A vssd1 vssd1 vccd1 vccd1 _13069_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10242_ _15497_/Q _10247_/C _10068_/X vssd1 vssd1 vccd1 vccd1 _10244_/C sky130_fd_sc_hd__a21o_1
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10173_ _10171_/B _10171_/C _10172_/X vssd1 vssd1 vccd1 vccd1 _10174_/C sky130_fd_sc_hd__o21ai_1
X_14981_ _16320_/Q _15131_/B _14981_/C vssd1 vssd1 vccd1 vccd1 _14984_/B sky130_fd_sc_hd__nand3_1
X_13932_ _13932_/A _13932_/B vssd1 vssd1 vccd1 vccd1 _16088_/D sky130_fd_sc_hd__nor2_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13863_ _14029_/A _13863_/B _13863_/C vssd1 vssd1 vccd1 vccd1 _13864_/A sky130_fd_sc_hd__and3_1
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15602_ _15602_/CLK _15602_/D vssd1 vssd1 vccd1 vccd1 _15602_/Q sky130_fd_sc_hd__dfxtp_2
X_12814_ _12813_/B _12813_/C _12758_/X vssd1 vssd1 vccd1 vccd1 _12815_/C sky130_fd_sc_hd__o21ai_1
X_13794_ _16067_/Q _13794_/B _13799_/C vssd1 vssd1 vccd1 vccd1 _13794_/Y sky130_fd_sc_hd__nand3_1
X_15533_ _15655_/CLK _15533_/D vssd1 vssd1 vccd1 vccd1 _15533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12745_ _12751_/A _12743_/Y _12744_/Y _12740_/C vssd1 vssd1 vccd1 vccd1 _12747_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _15484_/CLK _15464_/D vssd1 vssd1 vccd1 vccd1 _15464_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _15878_/Q _12684_/C _12616_/X vssd1 vssd1 vccd1 vccd1 _12676_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ _15014_/A vssd1 vssd1 vccd1 vccd1 _14415_/X sky130_fd_sc_hd__clkbuf_2
X_11627_ _11661_/A _11627_/B _11631_/A vssd1 vssd1 vccd1 vccd1 _15711_/D sky130_fd_sc_hd__nor3_1
X_15395_ _15395_/CLK _15395_/D vssd1 vssd1 vccd1 vccd1 _15395_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346_ _16176_/Q _14345_/C _14300_/X vssd1 vssd1 vccd1 vccd1 _14346_/Y sky130_fd_sc_hd__a21oi_1
X_11558_ _11597_/A _11558_/B _11558_/C vssd1 vssd1 vccd1 vccd1 _11559_/A sky130_fd_sc_hd__and3_1
XFILLER_7_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _10515_/A _10507_/Y _10508_/Y _10503_/C vssd1 vssd1 vccd1 vccd1 _10511_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14277_ _14321_/A _14277_/B vssd1 vssd1 vccd1 vccd1 _14277_/Y sky130_fd_sc_hd__nor2_1
X_11489_ _15691_/Q _11487_/C _11488_/X vssd1 vssd1 vccd1 vccd1 _11490_/B sky130_fd_sc_hd__a21oi_1
X_16016_ _16052_/CLK _16016_/D vssd1 vssd1 vccd1 vccd1 _16016_/Q sky130_fd_sc_hd__dfxtp_1
X_13228_ _13226_/X _13227_/Y _13222_/B _13223_/C vssd1 vssd1 vccd1 vccd1 _13230_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13172_/C vssd1 vssd1 vccd1 vccd1 _13187_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07720_ _16350_/Q vssd1 vssd1 vccd1 vccd1 _08127_/A sky130_fd_sc_hd__inv_2
XFILLER_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07651_ _07666_/A _07650_/Y _07638_/B _07639_/C vssd1 vssd1 vccd1 vccd1 _07653_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ _15354_/Q _09326_/C _09205_/X vssd1 vssd1 vccd1 vccd1 _09323_/C sky130_fd_sc_hd__a21o_1
X_09252_ _09251_/B _09251_/C _09019_/X vssd1 vssd1 vccd1 vccd1 _09253_/C sky130_fd_sc_hd__o21ai_1
X_08203_ _08203_/A _08082_/A vssd1 vssd1 vccd1 vccd1 _08203_/X sky130_fd_sc_hd__or2b_1
X_09183_ _09183_/A _09183_/B vssd1 vssd1 vccd1 vccd1 _09184_/B sky130_fd_sc_hd__nor2_1
X_08134_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08241_/B sky130_fd_sc_hd__xor2_4
X_08065_ _08065_/A vssd1 vssd1 vccd1 vccd1 _14627_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_134_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08967_ _08981_/C vssd1 vssd1 vccd1 vccd1 _08989_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07918_ _13523_/C _07918_/B vssd1 vssd1 vccd1 vccd1 _07952_/B sky130_fd_sc_hd__xnor2_2
X_08898_ _08897_/B _08897_/C _08726_/X vssd1 vssd1 vccd1 vccd1 _08899_/C sky130_fd_sc_hd__o21ai_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07849_ _10234_/A _07849_/B vssd1 vssd1 vccd1 vccd1 _07986_/A sky130_fd_sc_hd__xnor2_1
XFILLER_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _10916_/A _10863_/C vssd1 vssd1 vccd1 vccd1 _10860_/X sky130_fd_sc_hd__or2_1
XFILLER_25_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ _09519_/A _09519_/B _09519_/C vssd1 vssd1 vccd1 vccd1 _09520_/A sky130_fd_sc_hd__and3_1
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _11422_/A vssd1 vssd1 vccd1 vccd1 _11078_/B sky130_fd_sc_hd__buf_2
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12530_/A vssd1 vssd1 vccd1 vccd1 _15853_/D sky130_fd_sc_hd__clkbuf_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _12518_/A _12461_/B _12465_/B vssd1 vssd1 vccd1 vccd1 _15842_/D sky130_fd_sc_hd__nor3_1
XFILLER_149_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14200_ _14061_/X _14153_/X _14193_/B _13969_/X vssd1 vssd1 vccd1 vccd1 _14201_/B
+ sky130_fd_sc_hd__a31o_1
X_11412_ _11420_/A _11412_/B _11412_/C vssd1 vssd1 vccd1 vccd1 _11413_/A sky130_fd_sc_hd__and3_1
X_15180_ _15180_/A _15180_/B vssd1 vssd1 vccd1 vccd1 _15181_/B sky130_fd_sc_hd__nor2_1
XFILLER_137_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12392_ _15833_/Q _12399_/C _12332_/X vssd1 vssd1 vccd1 vccd1 _12392_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14131_ _16132_/Q _14137_/C _13893_/X vssd1 vssd1 vccd1 vccd1 _14133_/B sky130_fd_sc_hd__a21oi_1
X_11343_ _11343_/A _11343_/B _11343_/C vssd1 vssd1 vccd1 vccd1 _11344_/C sky130_fd_sc_hd__nand3_1
XFILLER_137_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ _14061_/X _15013_/A _14054_/B _13969_/X vssd1 vssd1 vccd1 vccd1 _14063_/B
+ sky130_fd_sc_hd__a31o_1
X_11274_ _15664_/Q _15663_/Q _15662_/Q _11273_/X vssd1 vssd1 vccd1 vccd1 _15656_/D
+ sky130_fd_sc_hd__o31a_1
X_13013_ _13011_/Y _13007_/C _13009_/X _13010_/Y vssd1 vssd1 vccd1 vccd1 _13014_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_134_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10225_ _10338_/A _10228_/C vssd1 vssd1 vccd1 vccd1 _10225_/X sky130_fd_sc_hd__or2_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10156_ _15483_/Q _10162_/C _09981_/X vssd1 vssd1 vccd1 vccd1 _10156_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _10085_/Y _10079_/C _10082_/X _10084_/Y vssd1 vssd1 vccd1 vccd1 _10088_/C
+ sky130_fd_sc_hd__a211o_1
X_14964_ _14964_/A vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13915_ _15005_/A vssd1 vssd1 vccd1 vccd1 _15186_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14895_ _14895_/A _14895_/B vssd1 vssd1 vccd1 vccd1 _16294_/D sky130_fd_sc_hd__nor2_1
XFILLER_35_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13846_ _16078_/Q _14093_/B _13846_/C vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__and3_1
X_13777_ _16065_/Q _14071_/B _13777_/C vssd1 vssd1 vccd1 vccd1 _13782_/A sky130_fd_sc_hd__and3_1
XFILLER_16_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10989_ _15613_/Q _11027_/C _10760_/X vssd1 vssd1 vccd1 vccd1 _10991_/B sky130_fd_sc_hd__a21oi_1
XFILLER_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15516_ _15655_/CLK _15516_/D vssd1 vssd1 vccd1 vccd1 _15516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12728_ _15886_/Q _12729_/C _12668_/X vssd1 vssd1 vccd1 vccd1 _12728_/Y sky130_fd_sc_hd__a21oi_1
X_15447_ _15484_/CLK _15447_/D vssd1 vssd1 vccd1 vccd1 _15447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ _12659_/A vssd1 vssd1 vccd1 vccd1 _15874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15378_ _15484_/CLK _15378_/D vssd1 vssd1 vccd1 vccd1 _15378_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ _14328_/X _14153_/X _14321_/B _14240_/X vssd1 vssd1 vccd1 vccd1 _14330_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _15437_/Q _10102_/B _09874_/C vssd1 vssd1 vccd1 vccd1 _09870_/Y sky130_fd_sc_hd__nand3_1
XFILLER_98_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08821_/A _08821_/B _08821_/C vssd1 vssd1 vccd1 vccd1 _08822_/A sky130_fd_sc_hd__and3_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08752_ _15266_/Q _08753_/C _08634_/X vssd1 vssd1 vccd1 vccd1 _08752_/Y sky130_fd_sc_hd__a21oi_1
X_07703_ _07703_/A _07703_/B vssd1 vssd1 vccd1 vccd1 _15204_/D sky130_fd_sc_hd__nor2_1
XFILLER_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08683_ _08704_/A _08683_/B _08683_/C vssd1 vssd1 vccd1 vccd1 _08684_/A sky130_fd_sc_hd__and3_1
X_07634_ _07634_/A vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__buf_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09304_ _10169_/A vssd1 vssd1 vccd1 vccd1 _09536_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09235_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__buf_2
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09166_ _13064_/B vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__buf_2
XFILLER_119_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08117_ _09367_/A _07728_/B _07727_/A vssd1 vssd1 vccd1 vccd1 _08242_/A sky130_fd_sc_hd__o21ai_4
X_09097_ _15319_/Q _09105_/C _08920_/X vssd1 vssd1 vccd1 vccd1 _09097_/Y sky130_fd_sc_hd__a21oi_1
X_08048_ _15827_/Q vssd1 vssd1 vccd1 vccd1 _12361_/A sky130_fd_sc_hd__inv_2
XFILLER_123_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10010_ _15461_/Q _10010_/B _10016_/C vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__nand3_1
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09999_ _10035_/A _09999_/B _09999_/C vssd1 vssd1 vccd1 vccd1 _10000_/A sky130_fd_sc_hd__and3_1
XFILLER_29_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11961_ _11961_/A vssd1 vssd1 vccd1 vccd1 _15763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10912_ _15601_/Q _10910_/C _10911_/X vssd1 vssd1 vccd1 vccd1 _10913_/B sky130_fd_sc_hd__a21oi_1
X_13700_ _13700_/A vssd1 vssd1 vccd1 vccd1 _14093_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14680_ _14680_/A _14680_/B vssd1 vssd1 vccd1 vccd1 _14682_/B sky130_fd_sc_hd__nor2_1
X_11892_ _15754_/Q _11891_/C _11775_/X vssd1 vssd1 vccd1 vccd1 _11893_/B sky130_fd_sc_hd__a21oi_1
X_13631_ _13631_/A _13631_/B _13631_/C vssd1 vssd1 vccd1 vccd1 _13632_/C sky130_fd_sc_hd__nand3_1
X_10843_ _10840_/X _10841_/Y _10842_/Y _10838_/C vssd1 vssd1 vccd1 vccd1 _10845_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16350_ _16352_/CLK _16350_/D vssd1 vssd1 vccd1 vccd1 _16350_/Q sky130_fd_sc_hd__dfxtp_1
X_13562_ _14653_/A vssd1 vssd1 vccd1 vccd1 _13562_/X sky130_fd_sc_hd__clkbuf_2
X_10774_ _10789_/A _10774_/B _10774_/C vssd1 vssd1 vccd1 vccd1 _10775_/A sky130_fd_sc_hd__and3_1
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15301_ _15301_/CLK _15301_/D vssd1 vssd1 vccd1 vccd1 _15301_/Q sky130_fd_sc_hd__dfxtp_1
X_12513_ _15852_/Q _12519_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12513_/Y sky130_fd_sc_hd__a21oi_1
X_16281_ _16283_/CLK _16281_/D vssd1 vssd1 vccd1 vccd1 _16281_/Q sky130_fd_sc_hd__dfxtp_2
X_13493_ _13490_/X _13491_/Y _13492_/Y _13488_/C vssd1 vssd1 vccd1 vccd1 _13495_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15232_ _15254_/CLK _15232_/D vssd1 vssd1 vccd1 vccd1 _15232_/Q sky130_fd_sc_hd__dfxtp_1
X_12444_ _12441_/X _12442_/Y _12443_/Y _12438_/C vssd1 vssd1 vccd1 vccd1 _12446_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ _16364_/Q _15163_/B _15165_/C vssd1 vssd1 vccd1 vccd1 _15168_/A sky130_fd_sc_hd__and3_1
XFILLER_138_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12375_ _12375_/A vssd1 vssd1 vccd1 vccd1 _15829_/D sky130_fd_sc_hd__clkbuf_1
X_14114_ _14117_/C vssd1 vssd1 vccd1 vccd1 _14125_/C sky130_fd_sc_hd__clkbuf_1
X_11326_ _11439_/A _11326_/B _11326_/C vssd1 vssd1 vccd1 vccd1 _11329_/B sky130_fd_sc_hd__or3_1
XFILLER_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15094_ _16346_/Q _15163_/B _15096_/C vssd1 vssd1 vccd1 vccd1 _15099_/A sky130_fd_sc_hd__and3_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14045_ _14041_/B _14040_/Y _14041_/A vssd1 vssd1 vccd1 vccd1 _14045_/Y sky130_fd_sc_hd__o21bai_1
X_11257_ _11255_/Y _11249_/C _11262_/A _11254_/Y vssd1 vssd1 vccd1 vccd1 _11262_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10208_ _10204_/X _10205_/Y _10207_/Y _10202_/C vssd1 vssd1 vccd1 vccd1 _10210_/B
+ sky130_fd_sc_hd__o211ai_1
X_11188_ _11186_/Y _11181_/C _11183_/X _11185_/Y vssd1 vssd1 vccd1 vccd1 _11189_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10139_ _10153_/A _10139_/B _10139_/C vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__and3_1
X_15996_ _16052_/CLK _15996_/D vssd1 vssd1 vccd1 vccd1 _15996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14947_ _14947_/A vssd1 vssd1 vccd1 vccd1 _16307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14878_ _14878_/A _14878_/B vssd1 vssd1 vccd1 vccd1 _14880_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13829_ _13829_/A _13829_/B _13829_/C vssd1 vssd1 vccd1 vccd1 _13830_/C sky130_fd_sc_hd__nand3_1
XFILLER_16_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ _09018_/B _09018_/C _09019_/X vssd1 vssd1 vccd1 vccd1 _09021_/C sky130_fd_sc_hd__o21ai_1
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09922_ _09922_/A _09922_/B _09922_/C vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__and3_1
XFILLER_113_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09853_ _15436_/Q _10022_/B _09855_/C vssd1 vssd1 vccd1 vccd1 _09853_/X sky130_fd_sc_hd__and3_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _08802_/X _08803_/Y _08799_/B _08800_/C vssd1 vssd1 vccd1 vccd1 _08806_/B
+ sky130_fd_sc_hd__o211ai_1
X_09784_ _15426_/Q _09784_/B _09784_/C vssd1 vssd1 vccd1 vccd1 _09784_/X sky130_fd_sc_hd__and3_1
XFILLER_105_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08735_ _08735_/A vssd1 vssd1 vccd1 vccd1 _08735_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08666_ _13972_/A vssd1 vssd1 vccd1 vccd1 _08704_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ input1/X vssd1 vssd1 vccd1 vccd1 _13043_/B sky130_fd_sc_hd__buf_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08597_ _13972_/A vssd1 vssd1 vccd1 vccd1 _08648_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09218_ _10081_/A vssd1 vssd1 vccd1 vccd1 _09444_/B sky130_fd_sc_hd__buf_2
X_10490_ _15535_/Q _10602_/B _10492_/C vssd1 vssd1 vccd1 vccd1 _10490_/X sky130_fd_sc_hd__and3_1
XFILLER_148_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09149_ _09149_/A _09149_/B _09149_/C vssd1 vssd1 vccd1 vccd1 _09150_/C sky130_fd_sc_hd__nand3_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _12157_/X _12158_/Y _12159_/Y _12154_/C vssd1 vssd1 vccd1 vccd1 _12162_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11111_ _11133_/A _11111_/B _11111_/C vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__and3_1
XFILLER_146_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12091_ _12091_/A vssd1 vssd1 vccd1 vccd1 _15784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11042_ _15628_/Q _15627_/Q _15626_/Q _10983_/X vssd1 vssd1 vccd1 vccd1 _15620_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15850_ _15907_/CLK _15850_/D vssd1 vssd1 vccd1 vccd1 _15850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14801_ _14799_/A _14799_/B _14800_/X vssd1 vssd1 vccd1 vccd1 _16273_/D sky130_fd_sc_hd__a21oi_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15781_ _15195_/Q _15781_/D vssd1 vssd1 vccd1 vccd1 _15781_/Q sky130_fd_sc_hd__dfxtp_1
X_12993_ _12993_/A _12993_/B _12993_/C vssd1 vssd1 vccd1 vccd1 _12994_/C sky130_fd_sc_hd__nand3_1
XFILLER_45_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14732_ _14694_/X _14730_/A _14695_/X vssd1 vssd1 vccd1 vccd1 _14733_/B sky130_fd_sc_hd__o21ai_1
X_11944_ _15762_/Q _11950_/C _11713_/X vssd1 vssd1 vccd1 vccd1 _11944_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11875_ _11883_/A _11875_/B _11875_/C vssd1 vssd1 vccd1 vccd1 _11876_/A sky130_fd_sc_hd__and3_1
X_14663_ _16247_/Q _14778_/B _14665_/C vssd1 vssd1 vccd1 vccd1 _14668_/A sky130_fd_sc_hd__and3_1
X_10826_ _15588_/Q _10835_/C _10655_/X vssd1 vssd1 vccd1 vccd1 _10826_/Y sky130_fd_sc_hd__a21oi_1
X_13614_ _13613_/B _13613_/C _13562_/X vssd1 vssd1 vccd1 vccd1 _13615_/C sky130_fd_sc_hd__o21ai_1
X_14594_ _16230_/Q _14593_/C _14634_/B vssd1 vssd1 vccd1 vccd1 _14594_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16333_ _16344_/CLK _16333_/D vssd1 vssd1 vccd1 vccd1 _16333_/Q sky130_fd_sc_hd__dfxtp_2
X_13545_ _13543_/Y _13538_/C _13541_/X _13542_/Y vssd1 vssd1 vccd1 vccd1 _13546_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10757_ _10770_/C vssd1 vssd1 vccd1 vccd1 _10778_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16264_ _16264_/CLK _16264_/D vssd1 vssd1 vccd1 vccd1 _16264_/Q sky130_fd_sc_hd__dfxtp_2
X_13476_ _13476_/A _13476_/B _13480_/A vssd1 vssd1 vccd1 vccd1 _16009_/D sky130_fd_sc_hd__nor3_1
X_10688_ _10688_/A _10688_/B vssd1 vssd1 vccd1 vccd1 _10690_/B sky130_fd_sc_hd__nor2_1
X_12427_ _12713_/A vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__clkbuf_4
X_15215_ _16304_/CLK _15215_/D vssd1 vssd1 vccd1 vccd1 state1[0] sky130_fd_sc_hd__dfxtp_2
X_16195_ _16204_/CLK _16195_/D vssd1 vssd1 vccd1 vccd1 _16195_/Q sky130_fd_sc_hd__dfxtp_1
X_15146_ _15146_/A _15146_/B vssd1 vssd1 vccd1 vccd1 _15147_/B sky130_fd_sc_hd__nor2_1
X_12358_ _12396_/A _12358_/B _12358_/C vssd1 vssd1 vccd1 vccd1 _12359_/A sky130_fd_sc_hd__and3_1
XFILLER_114_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ _11309_/A _11309_/B _11309_/C vssd1 vssd1 vccd1 vccd1 _11310_/A sky130_fd_sc_hd__and3_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15077_ _15181_/A _15077_/B vssd1 vssd1 vccd1 vccd1 _15077_/X sky130_fd_sc_hd__or2_1
X_12289_ _12287_/Y _12281_/C _12294_/A _12286_/Y vssd1 vssd1 vccd1 vccd1 _12294_/B
+ sky130_fd_sc_hd__a211oi_1
X_14028_ _14028_/A _14028_/B _14028_/C vssd1 vssd1 vccd1 vccd1 _14029_/C sky130_fd_sc_hd__nand3_1
XFILLER_95_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15979_ _15984_/CLK _15979_/D vssd1 vssd1 vccd1 vccd1 _15979_/Q sky130_fd_sc_hd__dfxtp_1
X_08520_ _08520_/A vssd1 vssd1 vccd1 vccd1 _15230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08451_ state1[6] vssd1 vssd1 vccd1 vccd1 _08453_/A sky130_fd_sc_hd__inv_2
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08382_ _08362_/A _08362_/B _08381_/Y vssd1 vssd1 vccd1 vccd1 _08389_/A sky130_fd_sc_hd__a21o_2
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09003_ _13598_/A vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_136_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09905_ _09903_/X _09904_/Y _09900_/B _09901_/C vssd1 vssd1 vccd1 vccd1 _09907_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09836_ _09867_/C vssd1 vssd1 vccd1 vccd1 _09874_/C sky130_fd_sc_hd__clkbuf_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09767_ _09767_/A vssd1 vssd1 vccd1 vccd1 _15421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _08718_/A _08718_/B vssd1 vssd1 vccd1 vccd1 _08719_/B sky130_fd_sc_hd__nor2_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _09775_/A _09698_/B _09703_/B vssd1 vssd1 vccd1 vccd1 _15410_/D sky130_fd_sc_hd__nor3_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08649_ _08649_/A vssd1 vssd1 vccd1 vccd1 _15248_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _11658_/Y _11653_/C _11665_/A _11656_/Y vssd1 vssd1 vccd1 vccd1 _11665_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _15554_/Q _10617_/C _10610_/X vssd1 vssd1 vccd1 vccd1 _10611_/Y sky130_fd_sc_hd__a21oi_1
X_11591_ _12734_/A vssd1 vssd1 vccd1 vccd1 _11819_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13330_ _13324_/B _13325_/C _13327_/X _13328_/Y vssd1 vssd1 vccd1 vccd1 _13331_/C
+ sky130_fd_sc_hd__a211o_1
X_10542_ _10540_/X _10541_/Y _10537_/B _10538_/C vssd1 vssd1 vccd1 vccd1 _10544_/B
+ sky130_fd_sc_hd__o211ai_1
X_13261_ _15987_/Q _15989_/Q _15988_/Q _13209_/X vssd1 vssd1 vccd1 vccd1 _15972_/D
+ sky130_fd_sc_hd__o31a_1
X_10473_ _13316_/A vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_108_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12212_ _12226_/A _12212_/B _12212_/C vssd1 vssd1 vccd1 vccd1 _12213_/A sky130_fd_sc_hd__and3_1
X_15000_ _14998_/A _14998_/B _14999_/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__a21oi_1
X_13192_ _13218_/A _13192_/B _13197_/B vssd1 vssd1 vccd1 vccd1 _15959_/D sky130_fd_sc_hd__nor3_1
X_12143_ _12713_/A vssd1 vssd1 vccd1 vccd1 _12369_/B sky130_fd_sc_hd__buf_2
XFILLER_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12074_ _12112_/A _12074_/B _12074_/C vssd1 vssd1 vccd1 vccd1 _12075_/A sky130_fd_sc_hd__and3_1
XFILLER_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11025_ _11023_/Y _11019_/C _11030_/A _11022_/Y vssd1 vssd1 vccd1 vccd1 _11030_/B
+ sky130_fd_sc_hd__a211oi_1
X_15902_ _07603_/A _15902_/D vssd1 vssd1 vccd1 vccd1 _15902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15833_ _15907_/CLK _15833_/D vssd1 vssd1 vccd1 vccd1 _15833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15764_ _15890_/CLK _15764_/D vssd1 vssd1 vccd1 vccd1 _15764_/Q sky130_fd_sc_hd__dfxtp_4
X_12976_ _12976_/A vssd1 vssd1 vccd1 vccd1 _13014_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14715_ _14709_/B _14710_/C _14721_/A _14713_/Y vssd1 vssd1 vccd1 vccd1 _14721_/B
+ sky130_fd_sc_hd__a211oi_1
X_11927_ _11941_/A _11927_/B _11927_/C vssd1 vssd1 vccd1 vccd1 _11928_/A sky130_fd_sc_hd__and3_1
X_15695_ _15794_/CLK _15695_/D vssd1 vssd1 vccd1 vccd1 _15695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14646_ _15043_/A vssd1 vssd1 vccd1 vccd1 _14646_/X sky130_fd_sc_hd__buf_2
XFILLER_21_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11858_ _15749_/Q _11863_/C _11798_/X vssd1 vssd1 vccd1 vccd1 _11860_/C sky130_fd_sc_hd__a21o_1
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10809_ _10809_/A vssd1 vssd1 vccd1 vccd1 _15583_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_19 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _15737_/Q vssd1 vssd1 vccd1 vccd1 _11804_/C sky130_fd_sc_hd__inv_2
X_14577_ _07701_/X _14573_/B _14814_/A vssd1 vssd1 vccd1 vccd1 _14579_/A sky130_fd_sc_hd__a21oi_1
X_16316_ _16317_/CLK _16316_/D vssd1 vssd1 vccd1 vccd1 _16316_/Q sky130_fd_sc_hd__dfxtp_2
X_13528_ _13529_/B _13529_/C _13529_/A vssd1 vssd1 vccd1 vccd1 _13530_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16247_ _16247_/CLK _16247_/D vssd1 vssd1 vccd1 vccd1 _16247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13459_ _15050_/A vssd1 vssd1 vccd1 vccd1 _13662_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16178_ _16187_/CLK _16178_/D vssd1 vssd1 vccd1 vccd1 _16178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15129_ _16355_/Q _15163_/B _15131_/C vssd1 vssd1 vccd1 vccd1 _15134_/A sky130_fd_sc_hd__and3_1
XFILLER_88_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07951_ _09658_/A _07892_/B _07891_/B vssd1 vssd1 vccd1 vccd1 _07984_/A sky130_fd_sc_hd__o21ai_2
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07882_ _07991_/A _07991_/B vssd1 vssd1 vccd1 vccd1 _07883_/B sky130_fd_sc_hd__xor2_4
XFILLER_95_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09621_ _15400_/Q _09733_/B _09623_/C vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__and3_1
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09552_ _09553_/B _09553_/C _09553_/A vssd1 vssd1 vccd1 vccd1 _09554_/B sky130_fd_sc_hd__a21o_1
X_08503_ _12661_/A vssd1 vssd1 vccd1 vccd1 _13534_/A sky130_fd_sc_hd__buf_6
XFILLER_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09483_ _09508_/C vssd1 vssd1 vccd1 vccd1 _09522_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08434_ state1[4] _08462_/B vssd1 vssd1 vccd1 vccd1 _08444_/B sky130_fd_sc_hd__and2_1
XFILLER_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08365_ _08365_/A vssd1 vssd1 vccd1 vccd1 _08365_/Y sky130_fd_sc_hd__inv_2
X_08296_ _08296_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__xnor2_4
XFILLER_20_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09819_ _09826_/B _09819_/B vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__or2_1
XFILLER_143_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12830_ _12851_/A _12830_/B _12830_/C vssd1 vssd1 vccd1 vccd1 _12831_/A sky130_fd_sc_hd__and3_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12761_/A vssd1 vssd1 vccd1 vccd1 _15889_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _16223_/Q _16222_/Q _16221_/Q _14421_/X vssd1 vssd1 vccd1 vccd1 _16206_/D
+ sky130_fd_sc_hd__o31a_1
X_11712_ _15726_/Q _11943_/B _11712_/C vssd1 vssd1 vccd1 vccd1 _11722_/A sky130_fd_sc_hd__and3_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _15483_/CLK _15480_/D vssd1 vssd1 vccd1 vccd1 _15480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12699_/B _12692_/B vssd1 vssd1 vccd1 vccd1 _12695_/A sky130_fd_sc_hd__or2_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _15714_/Q _11697_/B _11643_/C vssd1 vssd1 vccd1 vccd1 _11643_/Y sky130_fd_sc_hd__nand3_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14431_/A _14431_/B _14431_/C vssd1 vssd1 vccd1 vccd1 _14432_/C sky130_fd_sc_hd__nand3_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11574_ _11597_/A _11574_/B _11574_/C vssd1 vssd1 vccd1 vccd1 _11575_/A sky130_fd_sc_hd__and3_1
X_14362_ _14356_/Y _14357_/X _14359_/B vssd1 vssd1 vccd1 vccd1 _14365_/B sky130_fd_sc_hd__o21a_1
XFILLER_10_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16101_ _16119_/CLK _16101_/D vssd1 vssd1 vccd1 vccd1 _16101_/Q sky130_fd_sc_hd__dfxtp_2
X_10525_ _11963_/A vssd1 vssd1 vccd1 vccd1 _11099_/A sky130_fd_sc_hd__clkbuf_2
X_13313_ _13319_/C vssd1 vssd1 vccd1 vccd1 _13327_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14293_ _16166_/Q _14299_/C _14250_/X vssd1 vssd1 vccd1 vccd1 _14295_/C sky130_fd_sc_hd__a21o_1
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13244_ _13242_/Y _13237_/C _13249_/A _13241_/Y vssd1 vssd1 vccd1 vccd1 _13249_/B
+ sky130_fd_sc_hd__a211oi_1
X_16032_ _16040_/CLK _16032_/D vssd1 vssd1 vccd1 vccd1 _16032_/Q sky130_fd_sc_hd__dfxtp_1
X_10456_ _10456_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10457_/B sky130_fd_sc_hd__nor2_1
X_13175_ _13169_/B _13170_/C _13172_/X _13173_/Y vssd1 vssd1 vccd1 vccd1 _13176_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10387_ _10387_/A vssd1 vssd1 vccd1 vccd1 _15517_/D sky130_fd_sc_hd__clkbuf_1
X_12126_ _12126_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12130_/C sky130_fd_sc_hd__nor2_1
X_12057_ _15779_/Q _12174_/B _12062_/C vssd1 vssd1 vccd1 vccd1 _12057_/Y sky130_fd_sc_hd__nand3_1
XFILLER_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11008_ _15615_/Q _11121_/B _11008_/C vssd1 vssd1 vccd1 vccd1 _11008_/Y sky130_fd_sc_hd__nand3_1
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15816_ _15907_/CLK _15816_/D vssd1 vssd1 vccd1 vccd1 _15816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15747_ _15794_/CLK _15747_/D vssd1 vssd1 vccd1 vccd1 _15747_/Q sky130_fd_sc_hd__dfxtp_2
X_12959_ _12959_/A _12959_/B _12959_/C vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__and3_1
XFILLER_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ _15763_/CLK _15678_/D vssd1 vssd1 vccd1 vccd1 _15678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14629_ _14630_/B _14630_/C _14630_/A vssd1 vssd1 vccd1 vccd1 _14631_/B sky130_fd_sc_hd__a21o_1
X_08150_ _08264_/A _08264_/B vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__xor2_4
X_08081_ _08081_/A _08081_/B vssd1 vssd1 vccd1 vccd1 _08203_/A sky130_fd_sc_hd__xnor2_2
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08983_ _08981_/X _08982_/Y _08976_/B _08977_/C vssd1 vssd1 vccd1 vccd1 _08985_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_57_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ _09196_/A _07934_/B vssd1 vssd1 vccd1 vccd1 _07935_/B sky130_fd_sc_hd__xnor2_2
XFILLER_87_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ _15963_/Q _15981_/Q vssd1 vssd1 vccd1 vccd1 _08007_/B sky130_fd_sc_hd__xor2_2
XFILLER_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _09638_/C vssd1 vssd1 vccd1 vccd1 _09644_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_44_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07796_ _08065_/A _08066_/B vssd1 vssd1 vccd1 vccd1 _07797_/B sky130_fd_sc_hd__xnor2_2
X_09535_ _09533_/A _09533_/B _09534_/X vssd1 vssd1 vccd1 vccd1 _15384_/D sky130_fd_sc_hd__a21oi_1
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ _15376_/Q _09644_/B _09466_/C vssd1 vssd1 vccd1 vccd1 _09476_/B sky130_fd_sc_hd__and3_1
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08417_ hold16/X _15212_/Q _15211_/Q _07608_/X vssd1 vssd1 vccd1 vccd1 _15214_/D
+ sky130_fd_sc_hd__o31a_1
X_09397_ _15365_/Q _09403_/C _09166_/X vssd1 vssd1 vccd1 vccd1 _09397_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ _08349_/A _08349_/B _08349_/C vssd1 vssd1 vccd1 vccd1 _08386_/B sky130_fd_sc_hd__a21o_1
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08279_ _08279_/A vssd1 vssd1 vccd1 vccd1 _08403_/B sky130_fd_sc_hd__clkbuf_2
X_10310_ _15508_/Q _10310_/B _10312_/C vssd1 vssd1 vccd1 vccd1 _10310_/X sky130_fd_sc_hd__and3_1
X_11290_ _15660_/Q _11298_/C _11230_/X vssd1 vssd1 vccd1 vccd1 _11290_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10241_ _15497_/Q _10298_/B _10247_/C vssd1 vssd1 vccd1 vccd1 _10244_/B sky130_fd_sc_hd__nand3_1
X_10172_ _10751_/A vssd1 vssd1 vccd1 vccd1 _10172_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14980_ _14980_/A vssd1 vssd1 vccd1 vccd1 _15131_/B sky130_fd_sc_hd__clkbuf_2
X_13931_ _14413_/A _15013_/A _13917_/B _15184_/A vssd1 vssd1 vccd1 vccd1 _13932_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13862_ _13861_/B _13861_/C _13919_/A vssd1 vssd1 vccd1 vccd1 _13863_/C sky130_fd_sc_hd__o21ai_1
X_15601_ _15194_/Q _15601_/D vssd1 vssd1 vccd1 vccd1 _15601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12813_ _12869_/A _12813_/B _12813_/C vssd1 vssd1 vccd1 vccd1 _12815_/B sky130_fd_sc_hd__or3_1
XFILLER_62_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13793_ _16068_/Q _13799_/C _13693_/X vssd1 vssd1 vccd1 vccd1 _13793_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15532_ _15655_/CLK _15532_/D vssd1 vssd1 vccd1 vccd1 _15532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _15887_/Q _12744_/B _12748_/C vssd1 vssd1 vccd1 vccd1 _12744_/Y sky130_fd_sc_hd__nand3_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15483_/CLK _15463_/D vssd1 vssd1 vccd1 vccd1 _15463_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _15878_/Q _12675_/B _12684_/C vssd1 vssd1 vccd1 vccd1 _12675_/X sky130_fd_sc_hd__and3_1
X_14414_ _14414_/A vssd1 vssd1 vccd1 vccd1 _15014_/A sky130_fd_sc_hd__clkbuf_4
X_11626_ _15712_/Q _11737_/B _11635_/C vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__and3_1
X_15394_ _15484_/CLK _15394_/D vssd1 vssd1 vccd1 vccd1 _15394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14345_ _16176_/Q _14474_/B _14345_/C vssd1 vssd1 vccd1 vccd1 _14352_/A sky130_fd_sc_hd__and3_1
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11557_ _11556_/B _11556_/C _11327_/X vssd1 vssd1 vccd1 vccd1 _11558_/C sky130_fd_sc_hd__o21ai_1
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10508_ _15536_/Q _10681_/B _10512_/C vssd1 vssd1 vccd1 vccd1 _10508_/Y sky130_fd_sc_hd__nand3_1
XFILLER_144_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11488_ _11488_/A vssd1 vssd1 vccd1 vccd1 _11488_/X sky130_fd_sc_hd__clkbuf_2
X_14276_ _14320_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _14277_/B sky130_fd_sc_hd__and2_1
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16015_ _16022_/CLK _16015_/D vssd1 vssd1 vccd1 vccd1 _16015_/Q sky130_fd_sc_hd__dfxtp_1
X_10439_ _15527_/Q _10609_/B _10446_/C vssd1 vssd1 vccd1 vccd1 _10439_/X sky130_fd_sc_hd__and3_1
X_13227_ _15968_/Q _13226_/C _14869_/A vssd1 vssd1 vccd1 vccd1 _13227_/Y sky130_fd_sc_hd__a21oi_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _13162_/C vssd1 vssd1 vccd1 vccd1 _13172_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _15787_/Q _12223_/B _12115_/C vssd1 vssd1 vccd1 vccd1 _12109_/Y sky130_fd_sc_hd__nand3_1
X_13089_ _13089_/A vssd1 vssd1 vccd1 vccd1 _15944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07650_ _15204_/Q _07658_/C _07649_/X vssd1 vssd1 vccd1 vccd1 _07650_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09320_ _15354_/Q _09432_/B _09326_/C vssd1 vssd1 vccd1 vccd1 _09323_/B sky130_fd_sc_hd__nand3_1
XFILLER_81_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ _09419_/A _09251_/B _09251_/C vssd1 vssd1 vccd1 vccd1 _09253_/B sky130_fd_sc_hd__or3_1
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08202_ _08041_/A _08041_/B _08201_/Y vssd1 vssd1 vccd1 vccd1 _08221_/A sky130_fd_sc_hd__a21o_1
X_09182_ _09190_/B _09182_/B vssd1 vssd1 vccd1 vccd1 _09184_/A sky130_fd_sc_hd__or2_1
XFILLER_147_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08133_ _07740_/A _07740_/B _08132_/Y vssd1 vssd1 vccd1 vccd1 _08240_/B sky130_fd_sc_hd__o21a_1
XFILLER_119_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08064_ _08064_/A _08064_/B vssd1 vssd1 vccd1 vccd1 _08080_/A sky130_fd_sc_hd__xor2_4
XFILLER_108_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08966_ _08966_/A vssd1 vssd1 vccd1 vccd1 _08981_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07917_ _07960_/A _07917_/B vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__xnor2_4
X_08897_ _09133_/A _08897_/B _08897_/C vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__or3_1
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07848_ _11156_/A _07848_/B vssd1 vssd1 vccd1 vccd1 _07849_/B sky130_fd_sc_hd__xnor2_4
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07779_ _07779_/A _07779_/B vssd1 vssd1 vccd1 vccd1 _07780_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09518_ _09516_/Y _09511_/C _09514_/X _09515_/Y vssd1 vssd1 vccd1 vccd1 _09519_/C
+ sky130_fd_sc_hd__a211o_1
X_10790_ _10790_/A vssd1 vssd1 vccd1 vccd1 _15580_/D sky130_fd_sc_hd__clkbuf_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09458_/A _09449_/B _09449_/C vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__and3_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _12458_/Y _12454_/C _12465_/A _12457_/Y vssd1 vssd1 vccd1 vccd1 _12465_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_40_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11411_ _11409_/Y _11405_/C _11407_/X _11408_/Y vssd1 vssd1 vccd1 vccd1 _11412_/C
+ sky130_fd_sc_hd__a211o_1
X_12391_ _15833_/Q _12391_/B _12399_/C vssd1 vssd1 vccd1 vccd1 _12391_/X sky130_fd_sc_hd__and3_1
X_11342_ _11343_/B _11343_/C _11343_/A vssd1 vssd1 vccd1 vccd1 _11344_/B sky130_fd_sc_hd__a21o_1
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14130_ _16132_/Q _14221_/B _14137_/C vssd1 vssd1 vccd1 vccd1 _14133_/A sky130_fd_sc_hd__and3_1
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11273_ _12418_/A vssd1 vssd1 vccd1 vccd1 _11273_/X sky130_fd_sc_hd__buf_2
X_14061_ _14328_/A vssd1 vssd1 vccd1 vccd1 _14061_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10224_ _10224_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10228_/C sky130_fd_sc_hd__nor2_1
X_13012_ _13009_/X _13010_/Y _13011_/Y _13007_/C vssd1 vssd1 vccd1 vccd1 _13014_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10155_ _15483_/Q _10155_/B _10155_/C vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__and3_1
XFILLER_121_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10086_ _10082_/X _10084_/Y _10085_/Y _10079_/C vssd1 vssd1 vccd1 vccd1 _10088_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_58_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14963_ _14963_/A _14967_/C vssd1 vssd1 vccd1 vccd1 _14966_/A sky130_fd_sc_hd__and2_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_86_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15260_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13914_ _14363_/A vssd1 vssd1 vccd1 vccd1 _14054_/A sky130_fd_sc_hd__clkbuf_2
X_14894_ _14892_/X _14889_/A _14893_/X vssd1 vssd1 vccd1 vccd1 _14895_/B sky130_fd_sc_hd__o21ai_1
XFILLER_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _13845_/A vssd1 vssd1 vccd1 vccd1 _16075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13776_ _16065_/Q _13805_/C _13573_/X vssd1 vssd1 vccd1 vccd1 _13778_/B sky130_fd_sc_hd__a21oi_1
XFILLER_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10988_ _11021_/C vssd1 vssd1 vccd1 vccd1 _11027_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15515_ _15655_/CLK _15515_/D vssd1 vssd1 vccd1 vccd1 _15515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12727_ _15886_/Q _12947_/B _12729_/C vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__and3_1
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15446_ _15484_/CLK _15446_/D vssd1 vssd1 vccd1 vccd1 _15446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12658_ _12680_/A _12658_/B _12658_/C vssd1 vssd1 vccd1 vccd1 _12659_/A sky130_fd_sc_hd__and3_1
XFILLER_31_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11609_ _11609_/A _11609_/B vssd1 vssd1 vccd1 vccd1 _11614_/C sky130_fd_sc_hd__nor2_1
X_15377_ _15377_/CLK _15377_/D vssd1 vssd1 vccd1 vccd1 _15377_/Q sky130_fd_sc_hd__dfxtp_1
X_12589_ _12601_/C vssd1 vssd1 vccd1 vccd1 _12610_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_10_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _15845_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14328_ _14328_/A vssd1 vssd1 vccd1 vccd1 _14328_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14259_ _14253_/B _14254_/C _14264_/A _14257_/Y vssd1 vssd1 vccd1 vccd1 _14264_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_132_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ _08818_/Y _08814_/C _08816_/X _08817_/Y vssd1 vssd1 vccd1 vccd1 _08821_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _15266_/Q _08865_/B _08753_/C vssd1 vssd1 vccd1 vccd1 _08751_/X sky130_fd_sc_hd__and3_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15368_/CLK sky130_fd_sc_hd__clkbuf_16
X_07702_ _07701_/X _07692_/A _07690_/X vssd1 vssd1 vccd1 vccd1 _07703_/B sky130_fd_sc_hd__o21ai_1
X_08682_ _08682_/A _08682_/B _08682_/C vssd1 vssd1 vccd1 vccd1 _08683_/C sky130_fd_sc_hd__nand3_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07633_ _15203_/Q _14743_/B _07633_/C vssd1 vssd1 vccd1 vccd1 _07638_/B sky130_fd_sc_hd__nand3_1
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09303_ _09301_/A _09301_/B _09302_/X vssd1 vssd1 vccd1 vccd1 _15349_/D sky130_fd_sc_hd__a21oi_1
XFILLER_110_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09234_ _09234_/A vssd1 vssd1 vccd1 vccd1 _15338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09165_ _15330_/Q _09165_/B _09173_/C vssd1 vssd1 vccd1 vccd1 _09165_/X sky130_fd_sc_hd__and3_1
XFILLER_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08116_ _08116_/A _08236_/B vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__xnor2_4
XFILLER_119_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ _15319_/Q _09211_/B _09096_/C vssd1 vssd1 vccd1 vccd1 _09096_/X sky130_fd_sc_hd__and3_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08047_ _15809_/Q vssd1 vssd1 vccd1 vccd1 _12249_/A sky130_fd_sc_hd__inv_2
XFILLER_89_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09998_ _09997_/B _09997_/C _09884_/X vssd1 vssd1 vccd1 vccd1 _09999_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08949_ _08947_/Y _08942_/C _08954_/A _08946_/Y vssd1 vssd1 vccd1 vccd1 _08954_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_68_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15286_/CLK sky130_fd_sc_hd__clkbuf_16
X_11960_ _11997_/A _11960_/B _11960_/C vssd1 vssd1 vccd1 vccd1 _11961_/A sky130_fd_sc_hd__and3_1
XFILLER_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10911_ _11488_/A vssd1 vssd1 vccd1 vccd1 _10911_/X sky130_fd_sc_hd__buf_2
XFILLER_72_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11891_ _15754_/Q _12007_/B _11891_/C vssd1 vssd1 vccd1 vccd1 _11901_/B sky130_fd_sc_hd__and3_1
X_13630_ _13631_/B _13631_/C _13631_/A vssd1 vssd1 vccd1 vccd1 _13632_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10842_ _15589_/Q _11073_/B _10847_/C vssd1 vssd1 vccd1 vccd1 _10842_/Y sky130_fd_sc_hd__nand3_1
XFILLER_72_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ _13662_/A _13561_/B _13561_/C vssd1 vssd1 vccd1 vccd1 _13564_/B sky130_fd_sc_hd__or3_1
X_10773_ _10767_/B _10768_/C _10770_/X _10771_/Y vssd1 vssd1 vccd1 vccd1 _10774_/C
+ sky130_fd_sc_hd__a211o_1
X_15300_ _15312_/CLK _15300_/D vssd1 vssd1 vccd1 vccd1 _15300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12512_ _15852_/Q _12512_/B _12512_/C vssd1 vssd1 vccd1 vccd1 _12522_/A sky130_fd_sc_hd__and3_1
XFILLER_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16280_ _16283_/CLK _16280_/D vssd1 vssd1 vccd1 vccd1 _16280_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13492_ _16013_/Q _13543_/B _13498_/C vssd1 vssd1 vccd1 vccd1 _13492_/Y sky130_fd_sc_hd__nand3_1
XFILLER_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15231_ _15254_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 _15231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12443_ _15840_/Q _12554_/B _12443_/C vssd1 vssd1 vccd1 vccd1 _12443_/Y sky130_fd_sc_hd__nand3_1
XFILLER_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15162_ _16364_/Q _15176_/C _08735_/A vssd1 vssd1 vccd1 vccd1 _15164_/B sky130_fd_sc_hd__a21oi_1
X_12374_ _12396_/A _12374_/B _12374_/C vssd1 vssd1 vccd1 vccd1 _12375_/A sky130_fd_sc_hd__and3_1
X_14113_ _14434_/A vssd1 vssd1 vccd1 vccd1 _14208_/A sky130_fd_sc_hd__clkbuf_2
X_11325_ _11555_/A vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15093_ _16346_/Q _15107_/C _08735_/A vssd1 vssd1 vccd1 vccd1 _15095_/B sky130_fd_sc_hd__a21oi_1
XFILLER_141_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11256_ _11262_/A _11254_/Y _11255_/Y _11249_/C vssd1 vssd1 vccd1 vccd1 _11258_/B
+ sky130_fd_sc_hd__o211a_1
X_14044_ _14041_/A _14041_/B _14040_/Y _14043_/Y vssd1 vssd1 vccd1 vccd1 _16111_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_79_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10207_ _15490_/Q _10441_/B _10214_/C vssd1 vssd1 vccd1 vccd1 _10207_/Y sky130_fd_sc_hd__nand3_1
X_11187_ _11183_/X _11185_/Y _11186_/Y _11181_/C vssd1 vssd1 vccd1 vccd1 _11189_/B
+ sky130_fd_sc_hd__o211ai_1
X_10138_ _10131_/B _10132_/C _10135_/X _10136_/Y vssd1 vssd1 vccd1 vccd1 _10139_/C
+ sky130_fd_sc_hd__a211o_1
X_15995_ _16007_/CLK _15995_/D vssd1 vssd1 vccd1 vccd1 _15995_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_59_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _16337_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10069_ _15470_/Q _10074_/C _10068_/X vssd1 vssd1 vccd1 vccd1 _10071_/C sky130_fd_sc_hd__a21o_1
XFILLER_85_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14946_ _14946_/A _14946_/B _14946_/C vssd1 vssd1 vccd1 vccd1 _14947_/A sky130_fd_sc_hd__and3_1
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14877_ _14877_/A _14877_/B vssd1 vssd1 vccd1 vccd1 _14880_/A sky130_fd_sc_hd__or2_1
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13828_ _13829_/B _13829_/C _13829_/A vssd1 vssd1 vccd1 vccd1 _13830_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16368__17 vssd1 vssd1 vccd1 vccd1 _16368__17/HI io_oeb[0] sky130_fd_sc_hd__conb_1
X_13759_ _16061_/Q _13758_/C _13708_/X vssd1 vssd1 vccd1 vccd1 _13760_/B sky130_fd_sc_hd__a21oi_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15429_ _15484_/CLK _15429_/D vssd1 vssd1 vccd1 vccd1 _15429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09921_ _09919_/Y _09914_/C _09916_/X _09917_/Y vssd1 vssd1 vccd1 vccd1 _09922_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _09852_/A vssd1 vssd1 vccd1 vccd1 _15434_/D sky130_fd_sc_hd__clkbuf_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _15274_/Q _08811_/C _08625_/X vssd1 vssd1 vccd1 vccd1 _08803_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09783_/A vssd1 vssd1 vccd1 vccd1 _15424_/D sky130_fd_sc_hd__clkbuf_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08734_ _08769_/C vssd1 vssd1 vccd1 vccd1 _08775_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08665_ _08663_/A _08663_/B _08664_/X vssd1 vssd1 vccd1 vccd1 _15250_/D sky130_fd_sc_hd__a21oi_1
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _07633_/C vssd1 vssd1 vccd1 vccd1 _07658_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08596_ _08594_/A _08594_/B _08595_/X vssd1 vssd1 vccd1 vccd1 _15241_/D sky130_fd_sc_hd__a21oi_1
XFILLER_35_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09217_ _09217_/A vssd1 vssd1 vccd1 vccd1 _15336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09148_ _09149_/B _09149_/C _09149_/A vssd1 vssd1 vccd1 vccd1 _09150_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09079_ _15332_/Q _15331_/Q _15330_/Q _08901_/X vssd1 vssd1 vccd1 vccd1 _15315_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_135_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _11110_/A _11110_/B _11110_/C vssd1 vssd1 vccd1 vccd1 _11111_/C sky130_fd_sc_hd__nand3_1
X_12090_ _12112_/A _12090_/B _12090_/C vssd1 vssd1 vccd1 vccd1 _12091_/A sky130_fd_sc_hd__and3_1
XFILLER_122_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11041_ _11041_/A vssd1 vssd1 vccd1 vccd1 _15619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14800_ _14843_/A _14800_/B vssd1 vssd1 vccd1 vccd1 _14800_/X sky130_fd_sc_hd__or2_1
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15780_ _15195_/Q _15780_/D vssd1 vssd1 vccd1 vccd1 _15780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12992_ _12993_/B _12993_/C _12993_/A vssd1 vssd1 vccd1 vccd1 _12994_/B sky130_fd_sc_hd__a21o_1
XFILLER_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14731_ _14853_/A _14811_/B _14731_/C vssd1 vssd1 vccd1 vccd1 _14733_/A sky130_fd_sc_hd__and3_1
X_11943_ _15762_/Q _11943_/B _11943_/C vssd1 vssd1 vccd1 vccd1 _11953_/A sky130_fd_sc_hd__and3_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14662_ _16247_/Q _14677_/C _14503_/X vssd1 vssd1 vccd1 vccd1 _14664_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11874_ _11872_/Y _11867_/C _11870_/X _11871_/Y vssd1 vssd1 vccd1 vccd1 _11875_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13613_ _13662_/A _13613_/B _13613_/C vssd1 vssd1 vccd1 vccd1 _13615_/B sky130_fd_sc_hd__or3_1
X_10825_ _15588_/Q _10999_/B _10825_/C vssd1 vssd1 vccd1 vccd1 _10825_/X sky130_fd_sc_hd__and3_1
X_14593_ _16230_/Q _14593_/B _14593_/C vssd1 vssd1 vccd1 vccd1 _14600_/A sky130_fd_sc_hd__and3_1
X_16332_ _16352_/CLK _16332_/D vssd1 vssd1 vccd1 vccd1 _16332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13544_ _13541_/X _13542_/Y _13543_/Y _13538_/C vssd1 vssd1 vccd1 vccd1 _13546_/B
+ sky130_fd_sc_hd__o211ai_1
X_10756_ _15575_/Q vssd1 vssd1 vccd1 vccd1 _10770_/C sky130_fd_sc_hd__inv_2
XFILLER_41_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16263_ _16273_/CLK _16263_/D vssd1 vssd1 vccd1 vccd1 _16263_/Q sky130_fd_sc_hd__dfxtp_2
X_13475_ _16011_/Q _13675_/B _13475_/C vssd1 vssd1 vccd1 vccd1 _13480_/A sky130_fd_sc_hd__and3_1
X_10687_ _10694_/B _10687_/B vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__or2_1
X_15214_ _16353_/CLK _15214_/D vssd1 vssd1 vccd1 vccd1 spike_out[1] sky130_fd_sc_hd__dfxtp_4
X_12426_ _12518_/A _12426_/B _12431_/A vssd1 vssd1 vccd1 vccd1 _15837_/D sky130_fd_sc_hd__nor3_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16194_ _16204_/CLK _16194_/D vssd1 vssd1 vccd1 vccd1 _16194_/Q sky130_fd_sc_hd__dfxtp_1
X_15145_ _15145_/A _15145_/B vssd1 vssd1 vccd1 vccd1 _15146_/B sky130_fd_sc_hd__nor2_1
X_12357_ _12356_/B _12356_/C _12188_/X vssd1 vssd1 vccd1 vccd1 _12358_/C sky130_fd_sc_hd__o21ai_1
XFILLER_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11308_ _11306_/Y _11301_/C _11304_/X _11305_/Y vssd1 vssd1 vccd1 vccd1 _11309_/C
+ sky130_fd_sc_hd__a211o_1
X_15076_ _15076_/A _15076_/B vssd1 vssd1 vccd1 vccd1 _15077_/B sky130_fd_sc_hd__nor2_1
X_12288_ _12294_/A _12286_/Y _12287_/Y _12281_/C vssd1 vssd1 vccd1 vccd1 _12290_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14027_ _14028_/B _14028_/C _14028_/A vssd1 vssd1 vccd1 vccd1 _14029_/B sky130_fd_sc_hd__a21o_1
X_11239_ _15651_/Q _11409_/B _11239_/C vssd1 vssd1 vccd1 vccd1 _11239_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15978_ _16124_/CLK _15978_/D vssd1 vssd1 vccd1 vccd1 _15978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14929_ _14929_/A _14929_/B vssd1 vssd1 vccd1 vccd1 _16302_/D sky130_fd_sc_hd__nor2_1
XFILLER_24_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08450_ state1[6] _08462_/B _08452_/B vssd1 vssd1 vccd1 vccd1 _08465_/A sky130_fd_sc_hd__a21oi_2
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08381_ _08381_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _08381_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09002_ _15304_/Q _09008_/C _08824_/X vssd1 vssd1 vccd1 vccd1 _09002_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_145_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09904_ _15444_/Q _09911_/C _09786_/X vssd1 vssd1 vccd1 vccd1 _09904_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_116_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09835_ _09855_/C vssd1 vssd1 vccd1 vccd1 _09867_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09766_ _09807_/A _09766_/B _09766_/C vssd1 vssd1 vccd1 vccd1 _09767_/A sky130_fd_sc_hd__and3_1
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08717_ _08724_/B _08717_/B vssd1 vssd1 vccd1 vccd1 _08719_/A sky130_fd_sc_hd__or2_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09697_ _09695_/Y _09690_/C _09703_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _09703_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08648_ _08648_/A _08648_/B _08648_/C vssd1 vssd1 vccd1 vccd1 _08649_/A sky130_fd_sc_hd__and3_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _08577_/Y _08571_/C _08573_/X _08576_/Y vssd1 vssd1 vccd1 vccd1 _08580_/C
+ sky130_fd_sc_hd__a211o_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10610_/A vssd1 vssd1 vccd1 vccd1 _10610_/X sky130_fd_sc_hd__clkbuf_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11590_ input5/X vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10541_ _15543_/Q _10549_/C _10364_/X vssd1 vssd1 vccd1 vccd1 _10541_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _13153_/X _13257_/C _13259_/Y vssd1 vssd1 vccd1 vccd1 _15971_/D sky130_fd_sc_hd__a21oi_1
X_10472_ _10506_/C vssd1 vssd1 vccd1 vccd1 _10512_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_6_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12211_ _12204_/B _12205_/C _12208_/X _12209_/Y vssd1 vssd1 vccd1 vccd1 _12212_/C
+ sky130_fd_sc_hd__a211o_1
X_13191_ _13189_/Y _13184_/C _13197_/A _13188_/Y vssd1 vssd1 vccd1 vccd1 _13197_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _12234_/A _12142_/B _12147_/A vssd1 vssd1 vccd1 vccd1 _15792_/D sky130_fd_sc_hd__nor3_1
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12073_ _12072_/B _12072_/C _11902_/X vssd1 vssd1 vccd1 vccd1 _12074_/C sky130_fd_sc_hd__o21ai_1
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11024_ _11030_/A _11022_/Y _11023_/Y _11019_/C vssd1 vssd1 vccd1 vccd1 _11026_/B
+ sky130_fd_sc_hd__o211a_1
X_15901_ _07603_/A _15901_/D vssd1 vssd1 vccd1 vccd1 _15901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832_ _15907_/CLK _15832_/D vssd1 vssd1 vccd1 vccd1 _15832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15763_ _15763_/CLK _15763_/D vssd1 vssd1 vccd1 vccd1 _15763_/Q sky130_fd_sc_hd__dfxtp_1
X_12975_ _12973_/A _12973_/B _12974_/X vssd1 vssd1 vccd1 vccd1 _15924_/D sky130_fd_sc_hd__a21oi_1
XFILLER_17_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14714_ _14721_/A _14713_/Y _14709_/B _14710_/C vssd1 vssd1 vccd1 vccd1 _14716_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11926_ _11919_/B _11920_/C _11923_/X _11924_/Y vssd1 vssd1 vccd1 vccd1 _11927_/C
+ sky130_fd_sc_hd__a211o_1
X_15694_ _15794_/CLK _15694_/D vssd1 vssd1 vccd1 vccd1 _15694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14645_ _14643_/A _14643_/B _14644_/X vssd1 vssd1 vccd1 vccd1 _16237_/D sky130_fd_sc_hd__a21oi_1
X_11857_ _15749_/Q _12085_/B _11863_/C vssd1 vssd1 vccd1 vccd1 _11860_/B sky130_fd_sc_hd__nand3_1
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10808_ _10845_/A _10808_/B _10808_/C vssd1 vssd1 vccd1 vccd1 _10809_/A sky130_fd_sc_hd__and3_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14576_ _14413_/X _14573_/B _14575_/Y vssd1 vssd1 vccd1 vccd1 _16222_/D sky130_fd_sc_hd__o21a_1
X_11788_ _15745_/Q _15744_/Q _15743_/Q _11560_/X vssd1 vssd1 vccd1 vccd1 _15737_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16315_ _16317_/CLK _16315_/D vssd1 vssd1 vccd1 vccd1 _16315_/Q sky130_fd_sc_hd__dfxtp_2
X_13527_ _16021_/Q _13533_/C _13526_/X vssd1 vssd1 vccd1 vccd1 _13529_/C sky130_fd_sc_hd__a21o_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10739_ _10737_/Y _10732_/C _10744_/A _10735_/Y vssd1 vssd1 vccd1 vccd1 _10744_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_9_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16246_ _16247_/CLK _16246_/D vssd1 vssd1 vccd1 vccd1 _16246_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13458_ _13456_/A _13456_/B _13457_/X vssd1 vssd1 vccd1 vccd1 _16005_/D sky130_fd_sc_hd__a21oi_1
XFILLER_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12409_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__clkbuf_2
X_16177_ _16187_/CLK _16177_/D vssd1 vssd1 vccd1 vccd1 _16177_/Q sky130_fd_sc_hd__dfxtp_1
X_13389_ _15995_/Q _13543_/B _13394_/C vssd1 vssd1 vccd1 vccd1 _13389_/Y sky130_fd_sc_hd__nand3_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15128_ _16355_/Q _15142_/C _08735_/A vssd1 vssd1 vccd1 vccd1 _15130_/B sky130_fd_sc_hd__a21oi_1
XFILLER_141_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07950_ _07930_/A _07930_/B _07949_/X vssd1 vssd1 vccd1 vccd1 _08178_/A sky130_fd_sc_hd__o21a_2
X_15059_ _16337_/Q _15163_/B _15061_/C vssd1 vssd1 vccd1 vccd1 _15064_/A sky130_fd_sc_hd__and3_1
XFILLER_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07881_ _13937_/C _07881_/B vssd1 vssd1 vccd1 vccd1 _07991_/B sky130_fd_sc_hd__xnor2_2
XFILLER_96_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09620_ _09620_/A vssd1 vssd1 vccd1 vccd1 _15398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09551_ _15389_/Q _09557_/C _09490_/X vssd1 vssd1 vccd1 vccd1 _09553_/C sky130_fd_sc_hd__a21o_1
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08502_ _15230_/Q _08505_/C _12847_/A vssd1 vssd1 vccd1 vccd1 _08502_/Y sky130_fd_sc_hd__a21oi_1
X_09482_ _09496_/C vssd1 vssd1 vccd1 vccd1 _09508_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08433_ _08433_/A vssd1 vssd1 vccd1 vccd1 _08462_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08364_ _08391_/A _08391_/B vssd1 vssd1 vccd1 vccd1 _08368_/A sky130_fd_sc_hd__xor2_2
XFILLER_149_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08295_ _08295_/A _08295_/B vssd1 vssd1 vccd1 vccd1 _08296_/B sky130_fd_sc_hd__xnor2_2
XFILLER_133_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09818_ _15430_/Q _09817_/C _09755_/X vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__a21oi_1
XFILLER_74_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09749_ _15420_/Q _09754_/C _09693_/X vssd1 vssd1 vccd1 vccd1 _09749_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12796_/A _12760_/B _12760_/C vssd1 vssd1 vccd1 vccd1 _12761_/A sky130_fd_sc_hd__and3_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11711_ _12853_/A vssd1 vssd1 vccd1 vccd1 _11943_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _15880_/Q _12690_/C _12631_/X vssd1 vssd1 vccd1 vccd1 _12692_/B sky130_fd_sc_hd__a21oi_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14431_/B _14431_/C _14431_/A vssd1 vssd1 vccd1 vccd1 _14432_/B sky130_fd_sc_hd__a21o_1
X_11642_ _15715_/Q _11643_/C _11526_/X vssd1 vssd1 vccd1 vccd1 _11642_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _14356_/Y _14359_/X _14360_/Y vssd1 vssd1 vccd1 vccd1 _16175_/D sky130_fd_sc_hd__o21a_1
X_11573_ _11573_/A _11573_/B _11573_/C vssd1 vssd1 vccd1 vccd1 _11574_/C sky130_fd_sc_hd__nand3_1
XFILLER_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16100_ _16100_/CLK _16100_/D vssd1 vssd1 vccd1 vccd1 _16100_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13312_ _15972_/Q vssd1 vssd1 vccd1 vccd1 _13319_/C sky130_fd_sc_hd__inv_2
X_10524_ _15547_/Q _15546_/Q _15545_/Q _10409_/X vssd1 vssd1 vccd1 vccd1 _15539_/D
+ sky130_fd_sc_hd__o31a_1
X_14292_ _16166_/Q _14468_/B _14299_/C vssd1 vssd1 vccd1 vccd1 _14295_/B sky130_fd_sc_hd__nand3_1
X_16031_ _16031_/CLK _16031_/D vssd1 vssd1 vccd1 vccd1 _16031_/Q sky130_fd_sc_hd__dfxtp_1
X_13243_ _13249_/A _13241_/Y _13242_/Y _13237_/C vssd1 vssd1 vccd1 vccd1 _13245_/B
+ sky130_fd_sc_hd__o211a_1
X_10455_ _10463_/B _10455_/B vssd1 vssd1 vccd1 vccd1 _10457_/A sky130_fd_sc_hd__or2_1
XFILLER_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13174_ _13172_/X _13173_/Y _13169_/B _13170_/C vssd1 vssd1 vccd1 vccd1 _13176_/B
+ sky130_fd_sc_hd__o211ai_1
X_10386_ _10386_/A _10386_/B _10386_/C vssd1 vssd1 vccd1 vccd1 _10387_/A sky130_fd_sc_hd__and3_1
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12352_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _15780_/Q _12062_/C _12001_/X vssd1 vssd1 vccd1 vccd1 _12056_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _15616_/Q _11008_/C _10948_/X vssd1 vssd1 vccd1 vccd1 _11007_/Y sky130_fd_sc_hd__a21oi_1
X_15815_ _15907_/CLK _15815_/D vssd1 vssd1 vccd1 vccd1 _15815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15746_ _15746_/CLK _15746_/D vssd1 vssd1 vccd1 vccd1 _15746_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12958_ _12956_/Y _12952_/C _12954_/X _12955_/Y vssd1 vssd1 vccd1 vccd1 _12959_/C
+ sky130_fd_sc_hd__a211o_1
X_11909_ _11931_/C vssd1 vssd1 vccd1 vccd1 _11943_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15677_ _15763_/CLK _15677_/D vssd1 vssd1 vccd1 vccd1 _15677_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _12887_/X _12888_/Y _12884_/B _12885_/C vssd1 vssd1 vccd1 vccd1 _12891_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14628_ hold27/A _14627_/C _15165_/B vssd1 vssd1 vccd1 vccd1 _14630_/C sky130_fd_sc_hd__a21o_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14559_ _16222_/Q _14598_/B _14566_/C vssd1 vssd1 vccd1 vccd1 _14562_/A sky130_fd_sc_hd__and3_1
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _08080_/A _08080_/B vssd1 vssd1 vccd1 vccd1 _08081_/B sky130_fd_sc_hd__xor2_2
XFILLER_119_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16229_ _16362_/CLK _16229_/D vssd1 vssd1 vccd1 vccd1 _16229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08982_ _15301_/Q _08989_/C _08920_/X vssd1 vssd1 vccd1 vccd1 _08982_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07933_ _07933_/A _07933_/B vssd1 vssd1 vccd1 vccd1 _07934_/B sky130_fd_sc_hd__nand2_2
XFILLER_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07864_ _16116_/Q vssd1 vssd1 vccd1 vccd1 _14117_/C sky130_fd_sc_hd__inv_2
XFILLER_96_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09603_ _09623_/C vssd1 vssd1 vccd1 vccd1 _09638_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07795_ _15683_/Q _08072_/B vssd1 vssd1 vccd1 vccd1 _08066_/B sky130_fd_sc_hd__xnor2_4
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09534_ _09760_/A _09537_/C vssd1 vssd1 vccd1 vccd1 _09534_/X sky130_fd_sc_hd__or2_1
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09465_ _09487_/A _09465_/B _09470_/B vssd1 vssd1 vccd1 vccd1 _15374_/D sky130_fd_sc_hd__nor3_1
X_08416_ _08414_/X _08415_/Y _08412_/C _08471_/B vssd1 vssd1 vccd1 vccd1 _15213_/D
+ sky130_fd_sc_hd__a31oi_1
X_09396_ _15365_/Q _09451_/B _09403_/C vssd1 vssd1 vccd1 vccd1 _09396_/X sky130_fd_sc_hd__and3_1
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08347_ _08311_/A _08311_/B _08346_/Y vssd1 vssd1 vccd1 vccd1 _08349_/C sky130_fd_sc_hd__a21oi_1
XFILLER_138_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _08274_/Y _08276_/Y _08277_/Y vssd1 vssd1 vccd1 vccd1 _15208_/D sky130_fd_sc_hd__o21a_1
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10240_ _10353_/A _10240_/B _10244_/A vssd1 vssd1 vccd1 vccd1 _15495_/D sky130_fd_sc_hd__nor3_1
XFILLER_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10171_ _10284_/A _10171_/B _10171_/C vssd1 vssd1 vccd1 vccd1 _10174_/B sky130_fd_sc_hd__or3_1
XFILLER_78_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13930_ _13930_/A vssd1 vssd1 vccd1 vccd1 _15184_/A sky130_fd_sc_hd__buf_2
XFILLER_75_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13861_ _14106_/A _13861_/B _13861_/C vssd1 vssd1 vccd1 vccd1 _13863_/B sky130_fd_sc_hd__or3_1
XFILLER_28_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15600_ _15194_/Q _15600_/D vssd1 vssd1 vccd1 vccd1 _15600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12812_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12851_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13792_ _16068_/Q _13838_/B _13799_/C vssd1 vssd1 vccd1 vccd1 _13792_/X sky130_fd_sc_hd__and3_1
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15531_ _15655_/CLK _15531_/D vssd1 vssd1 vccd1 vccd1 _15531_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _15888_/Q _12748_/C _12569_/X vssd1 vssd1 vccd1 vccd1 _12743_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _15483_/CLK _15462_/D vssd1 vssd1 vccd1 vccd1 _15462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12674_/A vssd1 vssd1 vccd1 vccd1 _15876_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14413_/A vssd1 vssd1 vccd1 vccd1 _14413_/X sky130_fd_sc_hd__clkbuf_2
X_11625_ _15712_/Q _11662_/C _11624_/X vssd1 vssd1 vccd1 vccd1 _11627_/B sky130_fd_sc_hd__a21oi_1
X_15393_ _15484_/CLK _15393_/D vssd1 vssd1 vccd1 vccd1 _15393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14344_ _14344_/A vssd1 vssd1 vccd1 vccd1 _16172_/D sky130_fd_sc_hd__clkbuf_1
X_11556_ _11727_/A _11556_/B _11556_/C vssd1 vssd1 vccd1 vccd1 _11558_/B sky130_fd_sc_hd__or3_1
XFILLER_10_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10507_ _15537_/Q _10512_/C _10269_/X vssd1 vssd1 vccd1 vccd1 _10507_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14275_ _14268_/Y _14269_/X _14272_/B vssd1 vssd1 vccd1 vccd1 _14276_/B sky130_fd_sc_hd__o21a_1
X_11487_ _15691_/Q _11719_/B _11487_/C vssd1 vssd1 vccd1 vccd1 _11497_/B sky130_fd_sc_hd__and3_1
X_16014_ _16022_/CLK _16014_/D vssd1 vssd1 vccd1 vccd1 _16014_/Q sky130_fd_sc_hd__dfxtp_1
X_13226_ _15968_/Q _14298_/A _13226_/C vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__and3_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10438_ _10438_/A vssd1 vssd1 vccd1 vccd1 _15525_/D sky130_fd_sc_hd__clkbuf_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13157_ _15971_/Q _15970_/Q _15969_/Q _12981_/X vssd1 vssd1 vccd1 vccd1 _15954_/D
+ sky130_fd_sc_hd__o31a_1
X_10369_ _10369_/A vssd1 vssd1 vccd1 vccd1 _15515_/D sky130_fd_sc_hd__clkbuf_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _15788_/Q _12115_/C _12048_/X vssd1 vssd1 vccd1 vccd1 _12108_/Y sky130_fd_sc_hd__a21oi_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13088_ _13149_/A _13088_/B _13088_/C vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__and3_1
X_12039_ _15778_/Q _12099_/B _12042_/C vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__and3_1
XFILLER_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15729_ _15794_/CLK _15729_/D vssd1 vssd1 vccd1 vccd1 _15729_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09250_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09288_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08201_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08201_/Y sky130_fd_sc_hd__nor2_1
X_09181_ _15332_/Q _09179_/C _09180_/X vssd1 vssd1 vccd1 vccd1 _09182_/B sky130_fd_sc_hd__a21oi_1
X_08132_ _15972_/Q _08132_/B vssd1 vssd1 vccd1 vccd1 _08132_/Y sky130_fd_sc_hd__nand2_1
X_08063_ _08211_/B _08063_/B vssd1 vssd1 vccd1 vccd1 _08064_/B sky130_fd_sc_hd__nor2_2
XFILLER_147_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08965_ _15367_/Q _15366_/Q _15365_/Q _08901_/X vssd1 vssd1 vccd1 vccd1 _15297_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07916_ _07916_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07917_/B sky130_fd_sc_hd__nand2_2
XFILLER_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08896_ _11037_/A vssd1 vssd1 vccd1 vccd1 _09133_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07847_ _11275_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _07848_/B sky130_fd_sc_hd__xnor2_2
XFILLER_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07778_ _14706_/C _07778_/B vssd1 vssd1 vccd1 vccd1 _07779_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _09514_/X _09515_/Y _09516_/Y _09511_/C vssd1 vssd1 vccd1 vccd1 _09519_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09448_ _09446_/Y _09442_/C _09444_/X _09445_/Y vssd1 vssd1 vccd1 vccd1 _09449_/C
+ sky130_fd_sc_hd__a211o_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _09379_/A vssd1 vssd1 vccd1 vccd1 _15361_/D sky130_fd_sc_hd__clkbuf_1
X_11410_ _11407_/X _11408_/Y _11409_/Y _11405_/C vssd1 vssd1 vccd1 vccd1 _11412_/B
+ sky130_fd_sc_hd__o211ai_1
X_12390_ _12390_/A vssd1 vssd1 vccd1 vccd1 _15831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11341_ _15668_/Q _11347_/C _11222_/X vssd1 vssd1 vccd1 vccd1 _11343_/C sky130_fd_sc_hd__a21o_1
X_14060_ _14058_/X _14054_/B _14059_/X vssd1 vssd1 vccd1 vccd1 _14063_/A sky130_fd_sc_hd__a21oi_1
XFILLER_141_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11272_ _13720_/A vssd1 vssd1 vccd1 vccd1 _12418_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13011_ _15931_/Q _13066_/B _13016_/C vssd1 vssd1 vccd1 vccd1 _13011_/Y sky130_fd_sc_hd__nand3_1
X_10223_ _10223_/A _10223_/B vssd1 vssd1 vccd1 vccd1 _10224_/B sky130_fd_sc_hd__nor2_1
XFILLER_133_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10154_ _10154_/A vssd1 vssd1 vccd1 vccd1 _15481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14962_ _14802_/X _14955_/A _14958_/B _14961_/Y vssd1 vssd1 vccd1 vccd1 _16310_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_121_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10085_ _15471_/Q _10199_/B _10085_/C vssd1 vssd1 vccd1 vccd1 _10085_/Y sky130_fd_sc_hd__nand3_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13913_ _13901_/Y _13903_/X _13906_/B vssd1 vssd1 vccd1 vccd1 _13916_/B sky130_fd_sc_hd__o21a_1
X_14893_ _15169_/A vssd1 vssd1 vccd1 vccd1 _14893_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13844_ _13844_/A _13844_/B _13844_/C vssd1 vssd1 vccd1 vccd1 _13845_/A sky130_fd_sc_hd__and3_1
XFILLER_90_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13775_ _13799_/C vssd1 vssd1 vccd1 vccd1 _13805_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10987_ _11008_/C vssd1 vssd1 vccd1 vccd1 _11021_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15514_ _15655_/CLK _15514_/D vssd1 vssd1 vccd1 vccd1 _15514_/Q sky130_fd_sc_hd__dfxtp_1
X_12726_ _12726_/A vssd1 vssd1 vccd1 vccd1 _12947_/B sky130_fd_sc_hd__buf_2
XFILLER_30_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15445_ _15483_/CLK _15445_/D vssd1 vssd1 vccd1 vccd1 _15445_/Q sky130_fd_sc_hd__dfxtp_1
X_12657_ _12657_/A _12657_/B _12657_/C vssd1 vssd1 vccd1 vccd1 _12658_/C sky130_fd_sc_hd__nand3_1
XFILLER_129_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11608_ _11608_/A _11608_/B vssd1 vssd1 vccd1 vccd1 _11609_/B sky130_fd_sc_hd__nor2_1
X_15376_ _15484_/CLK _15376_/D vssd1 vssd1 vccd1 vccd1 _15376_/Q sky130_fd_sc_hd__dfxtp_1
X_12588_ _12588_/A vssd1 vssd1 vccd1 vccd1 _12601_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_117_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14327_ _14325_/X _14321_/B _14326_/X vssd1 vssd1 vccd1 vccd1 _14330_/A sky130_fd_sc_hd__a21oi_1
XFILLER_144_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11539_ _11539_/A vssd1 vssd1 vccd1 vccd1 _15697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14258_ _14264_/A _14257_/Y _14253_/B _14254_/C vssd1 vssd1 vccd1 vccd1 _14260_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13209_ _13723_/A vssd1 vssd1 vccd1 vccd1 _13209_/X sky130_fd_sc_hd__buf_2
XFILLER_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14183_/Y _14187_/X _14188_/Y vssd1 vssd1 vccd1 vccd1 _16139_/D sky130_fd_sc_hd__o21a_1
XFILLER_98_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08750_/A vssd1 vssd1 vccd1 vccd1 _15264_/D sky130_fd_sc_hd__clkbuf_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07701_ _14325_/A vssd1 vssd1 vccd1 vccd1 _07701_/X sky130_fd_sc_hd__buf_2
X_08681_ _08682_/B _08682_/C _08682_/A vssd1 vssd1 vccd1 vccd1 _08683_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ _07632_/A vssd1 vssd1 vccd1 vccd1 _14743_/B sky130_fd_sc_hd__buf_2
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09302_ _09472_/A _09306_/C vssd1 vssd1 vccd1 vccd1 _09302_/X sky130_fd_sc_hd__or2_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _09233_/A _09233_/B _09233_/C vssd1 vssd1 vccd1 vccd1 _09234_/A sky130_fd_sc_hd__and3_1
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09164_ _09164_/A vssd1 vssd1 vccd1 vccd1 _15328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08115_ _08115_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08236_/B sky130_fd_sc_hd__xor2_2
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09095_ _09095_/A vssd1 vssd1 vccd1 vccd1 _15317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08046_ _11502_/A _07785_/B _07784_/A vssd1 vssd1 vccd1 vccd1 _08081_/A sky130_fd_sc_hd__o21ai_2
XFILLER_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09997_ _09997_/A _09997_/B _09997_/C vssd1 vssd1 vccd1 vccd1 _09999_/B sky130_fd_sc_hd__or3_1
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08948_ _08954_/A _08946_/Y _08947_/Y _08942_/C vssd1 vssd1 vccd1 vccd1 _08950_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08879_ _08879_/A vssd1 vssd1 vccd1 vccd1 _15284_/D sky130_fd_sc_hd__clkbuf_1
X_10910_ _15601_/Q _11143_/B _10910_/C vssd1 vssd1 vccd1 vccd1 _10920_/B sky130_fd_sc_hd__and3_1
XFILLER_44_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11890_ _11949_/A _11890_/B _11894_/B vssd1 vssd1 vccd1 vccd1 _15752_/D sky130_fd_sc_hd__nor3_1
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _15590_/Q _10847_/C _10610_/X vssd1 vssd1 vccd1 vccd1 _10841_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ _13558_/A _13558_/B _13559_/X vssd1 vssd1 vccd1 vccd1 _16023_/D sky130_fd_sc_hd__a21oi_1
X_10772_ _10770_/X _10771_/Y _10767_/B _10768_/C vssd1 vssd1 vccd1 vccd1 _10774_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _12511_/A vssd1 vssd1 vccd1 vccd1 _15850_/D sky130_fd_sc_hd__clkbuf_1
X_13491_ _16014_/Q _13498_/C _13437_/X vssd1 vssd1 vccd1 vccd1 _13491_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15230_ _15230_/CLK _15230_/D vssd1 vssd1 vccd1 vccd1 _15230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ _15841_/Q _12443_/C _12384_/X vssd1 vssd1 vccd1 vccd1 _12442_/Y sky130_fd_sc_hd__a21oi_1
X_15161_ _15165_/C vssd1 vssd1 vccd1 vccd1 _15176_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12373_ _12373_/A _12373_/B _12373_/C vssd1 vssd1 vccd1 vccd1 _12374_/C sky130_fd_sc_hd__nand3_1
X_14112_ _16142_/Q _16141_/Q _16140_/Q _13973_/X vssd1 vssd1 vccd1 vccd1 _16125_/D
+ sky130_fd_sc_hd__o31a_1
X_11324_ _11612_/A vssd1 vssd1 vccd1 vccd1 _11555_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15092_ _15096_/C vssd1 vssd1 vccd1 vccd1 _15107_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14043_ _14041_/X _14040_/Y _14042_/X vssd1 vssd1 vccd1 vccd1 _14043_/Y sky130_fd_sc_hd__a21oi_1
X_11255_ _15653_/Q _11313_/B _11259_/C vssd1 vssd1 vccd1 vccd1 _11255_/Y sky130_fd_sc_hd__nand3_1
XFILLER_122_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ _10785_/A vssd1 vssd1 vccd1 vccd1 _10441_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_106_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11186_ _15643_/Q _11362_/B _11191_/C vssd1 vssd1 vccd1 vccd1 _11186_/Y sky130_fd_sc_hd__nand3_1
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10137_ _10135_/X _10136_/Y _10131_/B _10132_/C vssd1 vssd1 vccd1 vccd1 _10139_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15994_ _15994_/CLK _15994_/D vssd1 vssd1 vccd1 vccd1 _15994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10068_ _11222_/A vssd1 vssd1 vccd1 vccd1 _10068_/X sky130_fd_sc_hd__clkbuf_2
X_14945_ _14945_/A _14945_/B _14945_/C vssd1 vssd1 vccd1 vccd1 _14946_/C sky130_fd_sc_hd__nand3_1
XFILLER_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14876_ _16295_/Q _14875_/C _14718_/X vssd1 vssd1 vccd1 vccd1 _14877_/B sky130_fd_sc_hd__a21oi_1
XFILLER_63_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13827_ _16075_/Q _13832_/C _07634_/A vssd1 vssd1 vccd1 vccd1 _13829_/C sky130_fd_sc_hd__a21o_1
XFILLER_63_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13758_ _16061_/Q _13853_/B _13758_/C vssd1 vssd1 vccd1 vccd1 _13766_/B sky130_fd_sc_hd__and3_1
XFILLER_43_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12709_ _12742_/C vssd1 vssd1 vccd1 vccd1 _12748_/C sky130_fd_sc_hd__clkbuf_2
X_13689_ _13683_/B _13684_/C _13686_/X _13687_/Y vssd1 vssd1 vccd1 vccd1 _13690_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15428_ _15484_/CLK _15428_/D vssd1 vssd1 vccd1 vccd1 _15428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15359_ _15359_/CLK _15359_/D vssd1 vssd1 vccd1 vccd1 _15359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09920_ _09916_/X _09917_/Y _09919_/Y _09914_/C vssd1 vssd1 vccd1 vccd1 _09922_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09851_ _09865_/A _09851_/B _09851_/C vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__and3_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _15274_/Q _08919_/B _08802_/C vssd1 vssd1 vccd1 vccd1 _08802_/X sky130_fd_sc_hd__and3_1
XFILLER_85_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09807_/A _09782_/B _09782_/C vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__and3_1
XFILLER_39_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08753_/C vssd1 vssd1 vccd1 vccd1 _08769_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08893_/A _08667_/C vssd1 vssd1 vccd1 vccd1 _08664_/X sky130_fd_sc_hd__or2_1
XFILLER_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07615_ _07929_/A vssd1 vssd1 vccd1 vccd1 _07633_/C sky130_fd_sc_hd__buf_2
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08595_ _15030_/A _08600_/C vssd1 vssd1 vccd1 vccd1 _08595_/X sky130_fd_sc_hd__or2_1
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09216_ _09233_/A _09216_/B _09216_/C vssd1 vssd1 vccd1 vccd1 _09217_/A sky130_fd_sc_hd__and3_1
XFILLER_108_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09147_ _15327_/Q _09152_/C _08913_/X vssd1 vssd1 vccd1 vccd1 _09149_/C sky130_fd_sc_hd__a21o_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09078_ _09078_/A vssd1 vssd1 vccd1 vccd1 _15314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08029_ _15881_/Q vssd1 vssd1 vccd1 vccd1 _12706_/A sky130_fd_sc_hd__inv_2
X_11040_ _11076_/A _11040_/B _11040_/C vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__and3_1
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12991_ _15929_/Q _12996_/C _13099_/A vssd1 vssd1 vccd1 vccd1 _12993_/C sky130_fd_sc_hd__a21o_1
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11942_ _11942_/A vssd1 vssd1 vccd1 vccd1 _15760_/D sky130_fd_sc_hd__clkbuf_1
X_14730_ _14730_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _16257_/D sky130_fd_sc_hd__nor2_1
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14661_ _14665_/C vssd1 vssd1 vccd1 vccd1 _14677_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11873_ _11870_/X _11871_/Y _11872_/Y _11867_/C vssd1 vssd1 vccd1 vccd1 _11875_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13612_ _13612_/A vssd1 vssd1 vccd1 vccd1 _13664_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10824_ _10824_/A vssd1 vssd1 vccd1 vccd1 _15586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14592_ _14592_/A vssd1 vssd1 vccd1 vccd1 _16226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13543_ _16022_/Q _13543_/B _13548_/C vssd1 vssd1 vccd1 vccd1 _13543_/Y sky130_fd_sc_hd__nand3_1
X_16331_ _16337_/CLK _16331_/D vssd1 vssd1 vccd1 vccd1 _16331_/Q sky130_fd_sc_hd__dfxtp_1
X_10755_ _15583_/Q _15582_/Q _15581_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _15575_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16262_ _16273_/CLK _16262_/D vssd1 vssd1 vccd1 vccd1 _16262_/Q sky130_fd_sc_hd__dfxtp_2
X_13474_ _13474_/A vssd1 vssd1 vccd1 vccd1 _13675_/B sky130_fd_sc_hd__buf_2
X_10686_ _15565_/Q _10685_/C _10624_/X vssd1 vssd1 vccd1 vccd1 _10687_/B sky130_fd_sc_hd__a21oi_1
XFILLER_145_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15213_ _15254_/CLK _15213_/D vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dfxtp_1
X_12425_ _15838_/Q _12593_/B _12434_/C vssd1 vssd1 vccd1 vccd1 _12431_/A sky130_fd_sc_hd__and3_1
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16193_ _16204_/CLK _16193_/D vssd1 vssd1 vccd1 vccd1 _16193_/Q sky130_fd_sc_hd__dfxtp_1
X_15144_ _15144_/A _15144_/B vssd1 vssd1 vccd1 vccd1 _15146_/A sky130_fd_sc_hd__or2_1
X_12356_ _12583_/A _12356_/B _12356_/C vssd1 vssd1 vccd1 vccd1 _12358_/B sky130_fd_sc_hd__or3_1
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _11304_/X _11305_/Y _11306_/Y _11301_/C vssd1 vssd1 vccd1 vccd1 _11309_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15075_ _15075_/A _15075_/B vssd1 vssd1 vccd1 vccd1 _15076_/B sky130_fd_sc_hd__nor2_1
X_12287_ _15815_/Q _12458_/B _12291_/C vssd1 vssd1 vccd1 vccd1 _12287_/Y sky130_fd_sc_hd__nand3_1
XFILLER_113_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14026_ _16112_/Q _14032_/C _13982_/X vssd1 vssd1 vccd1 vccd1 _14028_/C sky130_fd_sc_hd__a21o_1
X_11238_ _15652_/Q _11239_/C _11237_/X vssd1 vssd1 vccd1 vccd1 _11238_/Y sky130_fd_sc_hd__a21oi_1
X_11169_ _15642_/Q _11289_/B _11169_/C vssd1 vssd1 vccd1 vccd1 _11169_/X sky130_fd_sc_hd__and3_1
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15977_ _16123_/CLK _15977_/D vssd1 vssd1 vccd1 vccd1 _15977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14928_ _14766_/X _14930_/C _14893_/X vssd1 vssd1 vccd1 vccd1 _14929_/B sky130_fd_sc_hd__o21ai_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14859_ _14863_/C vssd1 vssd1 vccd1 vccd1 _14875_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08380_ _08363_/B _08380_/B vssd1 vssd1 vccd1 vccd1 _08404_/A sky130_fd_sc_hd__and2b_2
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09001_ _15304_/Q _09001_/B _09001_/C vssd1 vssd1 vccd1 vccd1 _09011_/A sky130_fd_sc_hd__and3_1
XFILLER_145_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09903_ _15444_/Q _10074_/B _09903_/C vssd1 vssd1 vccd1 vccd1 _09903_/X sky130_fd_sc_hd__and3_1
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09834_ _09847_/C vssd1 vssd1 vccd1 vccd1 _09855_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09764_/B _09764_/C _09596_/X vssd1 vssd1 vccd1 vccd1 _09766_/C sky130_fd_sc_hd__o21ai_1
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08716_ _15260_/Q _08715_/C _08590_/X vssd1 vssd1 vccd1 vccd1 _08717_/B sky130_fd_sc_hd__a21oi_1
X_09696_ _09703_/A _09694_/Y _09695_/Y _09690_/C vssd1 vssd1 vccd1 vccd1 _09698_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08647_ _08645_/Y _08639_/C _08643_/X _08644_/Y vssd1 vssd1 vccd1 vccd1 _08648_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08578_ _08573_/X _08576_/Y _08577_/Y _08571_/C vssd1 vssd1 vccd1 vccd1 _08580_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10540_ _15543_/Q _10654_/B _10540_/C vssd1 vssd1 vccd1 vccd1 _10540_/X sky130_fd_sc_hd__and3_1
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ _10492_/C vssd1 vssd1 vccd1 vccd1 _10506_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12210_ _12208_/X _12209_/Y _12204_/B _12205_/C vssd1 vssd1 vccd1 vccd1 _12212_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_136_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13190_ _13197_/A _13188_/Y _13189_/Y _13184_/C vssd1 vssd1 vccd1 vccd1 _13192_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ _15793_/Q _12309_/B _12150_/C vssd1 vssd1 vccd1 vccd1 _12147_/A sky130_fd_sc_hd__and3_1
XFILLER_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ _12299_/A _12072_/B _12072_/C vssd1 vssd1 vccd1 vccd1 _12074_/B sky130_fd_sc_hd__or3_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11023_ _15617_/Q _11023_/B _11027_/C vssd1 vssd1 vccd1 vccd1 _11023_/Y sky130_fd_sc_hd__nand3_1
X_15900_ _07603_/A _15900_/D vssd1 vssd1 vccd1 vccd1 _15900_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15831_ _15907_/CLK _15831_/D vssd1 vssd1 vccd1 vccd1 _15831_/Q sky130_fd_sc_hd__dfxtp_1
X_15762_ _15763_/CLK _15762_/D vssd1 vssd1 vccd1 vccd1 _15762_/Q sky130_fd_sc_hd__dfxtp_1
X_12974_ _13199_/A _12977_/C vssd1 vssd1 vccd1 vccd1 _12974_/X sky130_fd_sc_hd__or2_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14713_ _16258_/Q _14717_/C _07649_/X vssd1 vssd1 vccd1 vccd1 _14713_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11925_ _11923_/X _11924_/Y _11919_/B _11920_/C vssd1 vssd1 vccd1 vccd1 _11927_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15693_ _15763_/CLK _15693_/D vssd1 vssd1 vccd1 vccd1 _15693_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11856_ _12713_/A vssd1 vssd1 vccd1 vccd1 _12085_/B sky130_fd_sc_hd__clkbuf_2
X_14644_ _14644_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14644_/X sky130_fd_sc_hd__or2_1
XFILLER_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10807_ _10806_/B _10806_/C _10751_/X vssd1 vssd1 vccd1 vccd1 _10808_/C sky130_fd_sc_hd__o21ai_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14575_ _13925_/X _14573_/B _14528_/X vssd1 vssd1 vccd1 vccd1 _14575_/Y sky130_fd_sc_hd__a21oi_1
X_11787_ _11787_/A vssd1 vssd1 vccd1 vccd1 _15736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16314_ _16344_/CLK _16314_/D vssd1 vssd1 vccd1 vccd1 _16314_/Q sky130_fd_sc_hd__dfxtp_1
X_13526_ _13526_/A vssd1 vssd1 vccd1 vccd1 _13526_/X sky130_fd_sc_hd__buf_2
X_10738_ _10744_/A _10735_/Y _10737_/Y _10732_/C vssd1 vssd1 vccd1 vccd1 _10740_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13457_ _13457_/A _13460_/C vssd1 vssd1 vccd1 vccd1 _13457_/X sky130_fd_sc_hd__or2_1
X_16245_ _16268_/CLK _16245_/D vssd1 vssd1 vccd1 vccd1 _16245_/Q sky130_fd_sc_hd__dfxtp_2
X_10669_ _10669_/A vssd1 vssd1 vccd1 vccd1 _15561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12408_ _12408_/A _12408_/B vssd1 vssd1 vccd1 vccd1 _12410_/B sky130_fd_sc_hd__nor2_1
X_13388_ _15996_/Q _13394_/C _13179_/X vssd1 vssd1 vccd1 vccd1 _13388_/Y sky130_fd_sc_hd__a21oi_1
X_16176_ _16187_/CLK _16176_/D vssd1 vssd1 vccd1 vccd1 _16176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15127_ _15131_/C vssd1 vssd1 vccd1 vccd1 _15142_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12339_ _15825_/Q _12512_/B _12339_/C vssd1 vssd1 vccd1 vccd1 _12350_/A sky130_fd_sc_hd__and3_1
XFILLER_126_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15058_ _16337_/Q _15072_/C _14901_/X vssd1 vssd1 vccd1 vccd1 _15060_/B sky130_fd_sc_hd__a21oi_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14009_ _14002_/Y _14003_/X _14006_/B vssd1 vssd1 vccd1 vccd1 _14010_/B sky130_fd_sc_hd__o21a_1
XFILLER_68_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07880_ _13777_/C _07880_/B vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__xnor2_4
XFILLER_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09550_ _15389_/Q _09721_/B _09557_/C vssd1 vssd1 vccd1 vccd1 _09553_/B sky130_fd_sc_hd__nand3_1
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08501_ _12668_/A vssd1 vssd1 vccd1 vccd1 _12847_/A sky130_fd_sc_hd__buf_2
X_09481_ _09481_/A vssd1 vssd1 vccd1 vccd1 _09496_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08432_ _08428_/Y _08430_/Y _08431_/Y vssd1 vssd1 vccd1 vccd1 _15217_/D sky130_fd_sc_hd__o21a_1
X_08363_ _08380_/B _08363_/B vssd1 vssd1 vccd1 vccd1 _08391_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08294_ _08207_/A _08207_/B _08209_/B _08209_/A vssd1 vssd1 vccd1 vccd1 _08295_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_149_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09817_ _15430_/Q _09931_/B _09817_/C vssd1 vssd1 vccd1 vccd1 _09826_/B sky130_fd_sc_hd__and3_1
XFILLER_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09748_ _15420_/Q _09867_/B _09748_/C vssd1 vssd1 vccd1 vccd1 _09758_/A sky130_fd_sc_hd__and3_1
XFILLER_100_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _10548_/A vssd1 vssd1 vccd1 vccd1 _09911_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11710_ input6/X vssd1 vssd1 vccd1 vccd1 _12853_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _15880_/Q _12861_/B _12690_/C vssd1 vssd1 vccd1 vccd1 _12699_/B sky130_fd_sc_hd__and3_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _15715_/Q _11811_/B _11643_/C vssd1 vssd1 vccd1 vccd1 _11641_/X sky130_fd_sc_hd__and3_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _14356_/Y _14359_/X _14316_/X vssd1 vssd1 vccd1 vccd1 _14360_/Y sky130_fd_sc_hd__a21oi_1
X_11572_ _11573_/B _11573_/C _11573_/A vssd1 vssd1 vccd1 vccd1 _11574_/B sky130_fd_sc_hd__a21o_1
XFILLER_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13311_ _15998_/Q _15997_/Q _15996_/Q _13209_/X vssd1 vssd1 vccd1 vccd1 _15981_/D
+ sky130_fd_sc_hd__o31a_1
X_10523_ _10523_/A vssd1 vssd1 vccd1 vccd1 _15538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14291_ _14291_/A vssd1 vssd1 vccd1 vccd1 _14468_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16030_ _16031_/CLK _16030_/D vssd1 vssd1 vccd1 vccd1 _16030_/Q sky130_fd_sc_hd__dfxtp_1
X_13242_ _15969_/Q _13293_/B _13246_/C vssd1 vssd1 vccd1 vccd1 _13242_/Y sky130_fd_sc_hd__nand3_1
X_10454_ _15529_/Q _10453_/C _10333_/X vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__a21oi_1
XFILLER_124_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ _15959_/Q _13172_/C _14869_/A vssd1 vssd1 vccd1 vccd1 _13173_/Y sky130_fd_sc_hd__a21oi_1
X_10385_ _10383_/Y _10378_/C _10381_/X _10382_/Y vssd1 vssd1 vccd1 vccd1 _10386_/C
+ sky130_fd_sc_hd__a211o_1
X_12124_ _12124_/A _12124_/B vssd1 vssd1 vccd1 vccd1 _12126_/B sky130_fd_sc_hd__nor2_1
XFILLER_111_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12055_ _15780_/Q _12228_/B _12055_/C vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__and3_1
XFILLER_78_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11006_ _15616_/Q _11236_/B _11008_/C vssd1 vssd1 vccd1 vccd1 _11006_/X sky130_fd_sc_hd__and3_1
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15814_ _07603_/A _15814_/D vssd1 vssd1 vccd1 vccd1 _15814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15745_ _15763_/CLK _15745_/D vssd1 vssd1 vccd1 vccd1 _15745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _12954_/X _12955_/Y _12956_/Y _12952_/C vssd1 vssd1 vccd1 vccd1 _12959_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11908_ _11923_/C vssd1 vssd1 vccd1 vccd1 _11931_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _15763_/CLK _15676_/D vssd1 vssd1 vccd1 vccd1 _15676_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _15912_/Q _12896_/C _12661_/X vssd1 vssd1 vccd1 vccd1 _12888_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14627_ hold27/A _14743_/B _14627_/C vssd1 vssd1 vccd1 vccd1 _14630_/B sky130_fd_sc_hd__nand3_1
X_11839_ _11839_/A _11839_/B vssd1 vssd1 vccd1 vccd1 _11843_/C sky130_fd_sc_hd__nor2_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14558_ _14626_/A _14558_/B _14561_/B vssd1 vssd1 vccd1 vccd1 _16218_/D sky130_fd_sc_hd__nor3_1
X_13509_ _13509_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13512_/C sky130_fd_sc_hd__nor2_1
XFILLER_146_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14489_ _14485_/Y _14488_/X _14415_/X vssd1 vssd1 vccd1 vccd1 _14489_/Y sky130_fd_sc_hd__a21oi_1
X_16228_ _16362_/CLK _16228_/D vssd1 vssd1 vccd1 vccd1 _16228_/Q sky130_fd_sc_hd__dfxtp_1
X_16159_ _16169_/CLK _16159_/D vssd1 vssd1 vccd1 vccd1 _16159_/Q sky130_fd_sc_hd__dfxtp_1
X_08981_ _15301_/Q _09211_/B _08981_/C vssd1 vssd1 vccd1 vccd1 _08981_/X sky130_fd_sc_hd__and3_1
XFILLER_130_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07932_ _15342_/Q _07932_/B vssd1 vssd1 vccd1 vccd1 _07933_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07863_ _16098_/Q vssd1 vssd1 vccd1 vccd1 _14022_/C sky130_fd_sc_hd__clkinv_2
X_09602_ _09615_/C vssd1 vssd1 vccd1 vccd1 _09623_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07794_ _15647_/Q _15665_/Q vssd1 vssd1 vccd1 vccd1 _08072_/B sky130_fd_sc_hd__xor2_4
XFILLER_56_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09533_ _09533_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _09537_/C sky130_fd_sc_hd__nor2_1
XFILLER_37_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09464_ _09462_/Y _09458_/C _09470_/A _09461_/Y vssd1 vssd1 vccd1 vccd1 _09470_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_52_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08415_ _08415_/A _08468_/A vssd1 vssd1 vccd1 vccd1 _08415_/Y sky130_fd_sc_hd__nand2_1
X_09395_ _09395_/A vssd1 vssd1 vccd1 vccd1 _15363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08346_ _08384_/B _08346_/B vssd1 vssd1 vccd1 vccd1 _08346_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_149_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08277_ _08274_/Y _08276_/Y _08168_/X vssd1 vssd1 vccd1 vccd1 _08277_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10170_ _10404_/A vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13860_ _14073_/A vssd1 vssd1 vccd1 vccd1 _14029_/A sky130_fd_sc_hd__buf_2
XFILLER_90_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12811_ _12809_/A _12809_/B _12810_/X vssd1 vssd1 vccd1 vccd1 _15897_/D sky130_fd_sc_hd__a21oi_1
XFILLER_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13791_ _14073_/A vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15530_ _15539_/CLK _15530_/D vssd1 vssd1 vccd1 vccd1 _15530_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _15888_/Q _12798_/B _12742_/C vssd1 vssd1 vccd1 vccd1 _12751_/A sky130_fd_sc_hd__and3_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _15483_/CLK _15461_/D vssd1 vssd1 vccd1 vccd1 _15461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12680_/A _12673_/B _12673_/C vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__and3_1
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11624_ _11624_/A vssd1 vssd1 vccd1 vccd1 _11624_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _14408_/X _14410_/B _14411_/Y vssd1 vssd1 vccd1 vccd1 _16185_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15392_ _15484_/CLK _15392_/D vssd1 vssd1 vccd1 vccd1 _15392_/Q sky130_fd_sc_hd__dfxtp_1
X_14343_ _14343_/A _14343_/B _14343_/C vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__and3_1
X_11555_ _11555_/A vssd1 vssd1 vccd1 vccd1 _11597_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10506_ _15537_/Q _10734_/B _10506_/C vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__and3_1
XFILLER_128_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14274_ _14268_/Y _14272_/X _14273_/Y vssd1 vssd1 vccd1 vccd1 _16157_/D sky130_fd_sc_hd__o21a_1
X_11486_ _12629_/A vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13225_ _13283_/A vssd1 vssd1 vccd1 vccd1 _13281_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16013_ _16022_/CLK _16013_/D vssd1 vssd1 vccd1 vccd1 _16013_/Q sky130_fd_sc_hd__dfxtp_1
X_10437_ _10444_/A _10437_/B _10437_/C vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__and3_1
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ _13153_/X _13149_/C _13155_/Y vssd1 vssd1 vccd1 vccd1 _15953_/D sky130_fd_sc_hd__a21oi_1
X_10368_ _10386_/A _10368_/B _10368_/C vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__and3_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _15788_/Q _12107_/B _12115_/C vssd1 vssd1 vccd1 vccd1 _12107_/X sky130_fd_sc_hd__and3_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13086_/B _13086_/C _14970_/A vssd1 vssd1 vccd1 vccd1 _13088_/C sky130_fd_sc_hd__o21ai_1
X_10299_ _15506_/Q _10304_/C _10068_/X vssd1 vssd1 vccd1 vccd1 _10301_/C sky130_fd_sc_hd__a21o_1
X_12038_ _12038_/A vssd1 vssd1 vccd1 vccd1 _15776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13989_ _14434_/A vssd1 vssd1 vccd1 vccd1 _14098_/A sky130_fd_sc_hd__clkbuf_2
X_15728_ _15728_/CLK _15728_/D vssd1 vssd1 vccd1 vccd1 _15728_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15659_ _15763_/CLK _15659_/D vssd1 vssd1 vccd1 vccd1 _15659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08200_ _08200_/A _08285_/A vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__xnor2_4
X_09180_ _10044_/A vssd1 vssd1 vccd1 vccd1 _09180_/X sky130_fd_sc_hd__buf_2
X_08131_ _08131_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__xnor2_4
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08062_ _08062_/A _08062_/B vssd1 vssd1 vccd1 vccd1 _08063_/B sky130_fd_sc_hd__and2_1
XFILLER_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08964_ _08964_/A vssd1 vssd1 vccd1 vccd1 _15296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07915_ hold28/A _16305_/Q vssd1 vssd1 vccd1 vccd1 _07916_/B sky130_fd_sc_hd__or2_1
XFILLER_124_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08895_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07846_ _12420_/A _07846_/B vssd1 vssd1 vccd1 vccd1 _08038_/B sky130_fd_sc_hd__xnor2_4
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07777_ _07777_/A vssd1 vssd1 vccd1 vccd1 _14706_/C sky130_fd_sc_hd__buf_6
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09516_ _15382_/Q _09572_/B _09522_/C vssd1 vssd1 vccd1 vccd1 _09516_/Y sky130_fd_sc_hd__nand3_1
XFILLER_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09447_ _09444_/X _09445_/Y _09446_/Y _09442_/C vssd1 vssd1 vccd1 vccd1 _09449_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09378_ _09401_/A _09378_/B _09378_/C vssd1 vssd1 vccd1 vccd1 _09379_/A sky130_fd_sc_hd__and3_1
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ _08329_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08330_/B sky130_fd_sc_hd__and2_1
XFILLER_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11340_ _15668_/Q _11510_/B _11347_/C vssd1 vssd1 vccd1 vccd1 _11343_/B sky130_fd_sc_hd__nand3_1
XFILLER_126_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ _11271_/A vssd1 vssd1 vccd1 vccd1 _15655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _15932_/Q _13016_/C _07672_/A vssd1 vssd1 vccd1 vccd1 _13010_/Y sky130_fd_sc_hd__a21oi_1
X_10222_ _10228_/B _10222_/B vssd1 vssd1 vccd1 vccd1 _10224_/A sky130_fd_sc_hd__or2_1
X_10153_ _10153_/A _10153_/B _10153_/C vssd1 vssd1 vccd1 vccd1 _10154_/A sky130_fd_sc_hd__and3_1
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10084_ _15472_/Q _10085_/C _10083_/X vssd1 vssd1 vccd1 vccd1 _10084_/Y sky130_fd_sc_hd__a21oi_1
X_14961_ _15045_/A _14967_/C vssd1 vssd1 vccd1 vccd1 _14961_/Y sky130_fd_sc_hd__nor2_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13912_ _14408_/A vssd1 vssd1 vccd1 vccd1 _13912_/X sky130_fd_sc_hd__clkbuf_2
X_14892_ _14892_/A vssd1 vssd1 vccd1 vccd1 _14892_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13843_ _13841_/Y _13836_/C _13838_/X _13839_/Y vssd1 vssd1 vccd1 vccd1 _13844_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13774_ _13785_/C vssd1 vssd1 vccd1 vccd1 _13799_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10986_ _10999_/C vssd1 vssd1 vccd1 vccd1 _11008_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15513_ _15655_/CLK _15513_/D vssd1 vssd1 vccd1 vccd1 _15513_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12725_ _12725_/A vssd1 vssd1 vccd1 vccd1 _15884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15444_ _15483_/CLK _15444_/D vssd1 vssd1 vccd1 vccd1 _15444_/Q sky130_fd_sc_hd__dfxtp_1
X_12656_ _12657_/B _12657_/C _12657_/A vssd1 vssd1 vccd1 vccd1 _12658_/B sky130_fd_sc_hd__a21o_1
XFILLER_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ _11614_/B _11607_/B vssd1 vssd1 vccd1 vccd1 _11609_/A sky130_fd_sc_hd__or2_1
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15375_ _15484_/CLK _15375_/D vssd1 vssd1 vccd1 vccd1 _15375_/Q sky130_fd_sc_hd__dfxtp_1
X_12587_ _15871_/Q _15870_/Q _15869_/Q _12418_/X vssd1 vssd1 vccd1 vccd1 _15863_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_129_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14326_ _14326_/A vssd1 vssd1 vccd1 vccd1 _14326_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11538_ _11538_/A _11538_/B _11538_/C vssd1 vssd1 vccd1 vccd1 _11539_/A sky130_fd_sc_hd__and3_1
XFILLER_129_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14257_ _16158_/Q _14256_/C _14033_/X vssd1 vssd1 vccd1 vccd1 _14257_/Y sky130_fd_sc_hd__a21oi_1
X_11469_ _11477_/A _11469_/B _11469_/C vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__and3_1
XFILLER_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13208_ _13153_/X _13204_/C _13207_/Y vssd1 vssd1 vccd1 vccd1 _15962_/D sky130_fd_sc_hd__a21oi_1
X_14188_ _14183_/Y _14187_/X _14049_/X vssd1 vssd1 vccd1 vccd1 _14188_/Y sky130_fd_sc_hd__a21oi_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13139_ _15953_/Q _13138_/C _14364_/A vssd1 vssd1 vccd1 vccd1 _13140_/B sky130_fd_sc_hd__a21oi_1
XFILLER_124_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07700_ _14653_/A vssd1 vssd1 vccd1 vccd1 _14325_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08680_ _15255_/Q _08686_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _08682_/C sky130_fd_sc_hd__a21o_1
XFILLER_66_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07631_ _07634_/A vssd1 vssd1 vccd1 vccd1 _07632_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ _09301_/A _09301_/B vssd1 vssd1 vccd1 vccd1 _09306_/C sky130_fd_sc_hd__nor2_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ _09230_/Y _09225_/C _09228_/X _09229_/Y vssd1 vssd1 vccd1 vccd1 _09233_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09163_ _09171_/A _09163_/B _09163_/C vssd1 vssd1 vccd1 vccd1 _09164_/A sky130_fd_sc_hd__and3_1
XFILLER_147_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08114_ _09601_/A _09481_/A _08113_/Y vssd1 vssd1 vccd1 vccd1 _08115_/B sky130_fd_sc_hd__o21ai_4
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09094_ _09115_/A _09094_/B _09094_/C vssd1 vssd1 vccd1 vccd1 _09095_/A sky130_fd_sc_hd__and3_1
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08045_ _11388_/A _07800_/B _08044_/X vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__o21ai_4
XFILLER_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09996_ _10114_/A vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08947_ _15294_/Q _08947_/B _08951_/C vssd1 vssd1 vccd1 vccd1 _08947_/Y sky130_fd_sc_hd__nand3_1
XFILLER_57_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08878_ _08878_/A _08878_/B _08878_/C vssd1 vssd1 vccd1 vccd1 _08879_/A sky130_fd_sc_hd__and3_1
XFILLER_45_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07829_ _15368_/Q _08148_/B vssd1 vssd1 vccd1 vccd1 _07893_/A sky130_fd_sc_hd__xnor2_4
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10840_ _15590_/Q _10895_/B _10847_/C vssd1 vssd1 vccd1 vccd1 _10840_/X sky130_fd_sc_hd__and3_1
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ _15579_/Q _10778_/C _10655_/X vssd1 vssd1 vccd1 vccd1 _10771_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12510_ _12510_/A _12510_/B _12510_/C vssd1 vssd1 vccd1 vccd1 _12511_/A sky130_fd_sc_hd__and3_1
XFILLER_13_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13490_ _16014_/Q _13589_/B _13498_/C vssd1 vssd1 vccd1 vccd1 _13490_/X sky130_fd_sc_hd__and3_1
XFILLER_9_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12441_ _15841_/Q _12667_/B _12443_/C vssd1 vssd1 vccd1 vccd1 _12441_/X sky130_fd_sc_hd__and3_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12372_ _12373_/B _12373_/C _12373_/A vssd1 vssd1 vccd1 vccd1 _12374_/B sky130_fd_sc_hd__a21o_1
X_15160_ _15205_/Q _15204_/Q _15203_/Q _15017_/X vssd1 vssd1 vccd1 vccd1 _16359_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11323_ _11321_/A _11321_/B _11322_/X vssd1 vssd1 vccd1 vccd1 _15663_/D sky130_fd_sc_hd__a21oi_1
X_14111_ _13154_/X _14108_/C _14110_/Y vssd1 vssd1 vccd1 vccd1 _16124_/D sky130_fd_sc_hd__a21oi_1
X_15091_ _16358_/Q _16357_/Q _16356_/Q _15017_/X vssd1 vssd1 vccd1 vccd1 _16341_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11254_ _15654_/Q _11259_/C _11137_/X vssd1 vssd1 vccd1 vccd1 _11254_/Y sky130_fd_sc_hd__a21oi_1
X_14042_ _14883_/A vssd1 vssd1 vccd1 vccd1 _14042_/X sky130_fd_sc_hd__buf_2
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _15491_/Q _10214_/C _10030_/X vssd1 vssd1 vccd1 vccd1 _10205_/Y sky130_fd_sc_hd__a21oi_1
X_11185_ _15644_/Q _11191_/C _11184_/X vssd1 vssd1 vccd1 vccd1 _11185_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ _15480_/Q _10143_/C _10075_/X vssd1 vssd1 vccd1 vccd1 _10136_/Y sky130_fd_sc_hd__a21oi_1
X_15993_ _16007_/CLK _15993_/D vssd1 vssd1 vccd1 vccd1 _15993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10067_ input2/X vssd1 vssd1 vccd1 vccd1 _11222_/A sky130_fd_sc_hd__buf_4
X_14944_ _14945_/B _14945_/C _14945_/A vssd1 vssd1 vccd1 vccd1 _14946_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14875_ _16295_/Q _14953_/B _14875_/C vssd1 vssd1 vccd1 vccd1 _14877_/A sky130_fd_sc_hd__and3_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13826_ _16075_/Q _14074_/B _13832_/C vssd1 vssd1 vccd1 vccd1 _13829_/B sky130_fd_sc_hd__nand3_1
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ _13852_/A _13757_/B _13761_/B vssd1 vssd1 vccd1 vccd1 _16058_/D sky130_fd_sc_hd__nor3_1
X_10969_ _10969_/A vssd1 vssd1 vccd1 vccd1 _10970_/C sky130_fd_sc_hd__buf_2
X_12708_ _12729_/C vssd1 vssd1 vccd1 vccd1 _12742_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13688_ _13686_/X _13687_/Y _13683_/B _13684_/C vssd1 vssd1 vccd1 vccd1 _13690_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_31_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15427_ _15483_/CLK _15427_/D vssd1 vssd1 vccd1 vccd1 _15427_/Q sky130_fd_sc_hd__dfxtp_1
X_12639_ _12639_/A vssd1 vssd1 vccd1 vccd1 _12869_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15358_ _15359_/CLK _15358_/D vssd1 vssd1 vccd1 vccd1 _15358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14309_ _14883_/A vssd1 vssd1 vccd1 vccd1 _14309_/X sky130_fd_sc_hd__buf_2
X_15289_ _16344_/CLK _15289_/D vssd1 vssd1 vccd1 vccd1 _15289_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09850_ _09843_/B _09844_/C _09847_/X _09848_/Y vssd1 vssd1 vccd1 vccd1 _09851_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08801_ _08801_/A vssd1 vssd1 vccd1 vccd1 _15272_/D sky130_fd_sc_hd__clkbuf_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09781_/A _09781_/B _09781_/C vssd1 vssd1 vccd1 vccd1 _09782_/C sky130_fd_sc_hd__nand3_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _08745_/C vssd1 vssd1 vccd1 vccd1 _08753_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08663_ _08663_/A _08663_/B vssd1 vssd1 vccd1 vccd1 _08667_/C sky130_fd_sc_hd__nor2_1
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07614_ _16359_/Q vssd1 vssd1 vccd1 vccd1 _07929_/A sky130_fd_sc_hd__inv_2
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08594_ _08594_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08600_/C sky130_fd_sc_hd__nor2_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09215_ _09208_/B _09209_/C _09211_/X _09213_/Y vssd1 vssd1 vccd1 vccd1 _09216_/C
+ sky130_fd_sc_hd__a211o_1
X_09146_ _15327_/Q _09146_/B _09152_/C vssd1 vssd1 vccd1 vccd1 _09149_/B sky130_fd_sc_hd__nand3_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09077_ _09115_/A _09077_/B _09077_/C vssd1 vssd1 vccd1 vccd1 _09078_/A sky130_fd_sc_hd__and3_1
XFILLER_107_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08028_ _15863_/Q vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__inv_2
XFILLER_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09979_ _15456_/Q _10155_/B _09979_/C vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__and3_1
XFILLER_130_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12990_ _15929_/Q _13045_/B _12996_/C vssd1 vssd1 vccd1 vccd1 _12993_/B sky130_fd_sc_hd__nand3_1
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11941_ _11941_/A _11941_/B _11941_/C vssd1 vssd1 vccd1 vccd1 _11942_/A sky130_fd_sc_hd__and3_1
X_14660_ _16233_/Q vssd1 vssd1 vccd1 vccd1 _14665_/C sky130_fd_sc_hd__inv_2
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11872_ _15750_/Q _11986_/B _11872_/C vssd1 vssd1 vccd1 vccd1 _11872_/Y sky130_fd_sc_hd__nand3_1
XFILLER_60_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13611_ _13609_/A _13609_/B _13610_/X vssd1 vssd1 vccd1 vccd1 _16032_/D sky130_fd_sc_hd__a21oi_1
X_10823_ _10845_/A _10823_/B _10823_/C vssd1 vssd1 vccd1 vccd1 _10824_/A sky130_fd_sc_hd__and3_1
X_14591_ _14748_/A _14591_/B _14591_/C vssd1 vssd1 vccd1 vccd1 _14592_/A sky130_fd_sc_hd__and3_1
X_16330_ _16337_/CLK _16330_/D vssd1 vssd1 vccd1 vccd1 _16330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13542_ _16023_/Q _13548_/C _13437_/X vssd1 vssd1 vccd1 vccd1 _13542_/Y sky130_fd_sc_hd__a21oi_1
X_10754_ _10754_/A vssd1 vssd1 vccd1 vccd1 _15574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _16273_/CLK _16261_/D vssd1 vssd1 vccd1 vccd1 _16261_/Q sky130_fd_sc_hd__dfxtp_2
X_10685_ _15565_/Q _10798_/B _10685_/C vssd1 vssd1 vccd1 vccd1 _10694_/B sky130_fd_sc_hd__and3_1
XFILLER_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13473_ _16011_/Q _13504_/C _13317_/X vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__a21oi_1
X_15212_ _16224_/CLK _15212_/D vssd1 vssd1 vccd1 vccd1 _15212_/Q sky130_fd_sc_hd__dfxtp_1
X_16373__22 vssd1 vssd1 vccd1 vccd1 _16373__22/HI io_oeb[5] sky130_fd_sc_hd__conb_1
X_12424_ _15838_/Q _12462_/C _12197_/X vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__a21oi_1
X_16192_ _16192_/CLK _16192_/D vssd1 vssd1 vccd1 vccd1 _16192_/Q sky130_fd_sc_hd__dfxtp_1
X_15143_ _16358_/Q _15142_/C _13950_/B vssd1 vssd1 vccd1 vccd1 _15144_/B sky130_fd_sc_hd__a21oi_1
X_12355_ _12639_/A vssd1 vssd1 vccd1 vccd1 _12583_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ _15661_/Q _11362_/B _11311_/C vssd1 vssd1 vccd1 vccd1 _11306_/Y sky130_fd_sc_hd__nand3_1
X_12286_ _15816_/Q _12291_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12286_/Y sky130_fd_sc_hd__a21oi_1
X_15074_ _15074_/A _15074_/B vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__or2_1
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11237_ _12100_/A vssd1 vssd1 vccd1 vccd1 _11237_/X sky130_fd_sc_hd__buf_2
X_14025_ _16112_/Q _14249_/B _14032_/C vssd1 vssd1 vccd1 vccd1 _14028_/B sky130_fd_sc_hd__nand3_1
XFILLER_106_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11168_ _11168_/A vssd1 vssd1 vccd1 vccd1 _15640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10119_ _10983_/A vssd1 vssd1 vccd1 vccd1 _10119_/X sky130_fd_sc_hd__clkbuf_2
X_11099_ _11099_/A vssd1 vssd1 vccd1 vccd1 _11220_/A sky130_fd_sc_hd__buf_2
XFILLER_110_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15976_ _15984_/CLK _15976_/D vssd1 vssd1 vccd1 vccd1 _15976_/Q sky130_fd_sc_hd__dfxtp_1
X_14927_ _14963_/A _14930_/C vssd1 vssd1 vccd1 vccd1 _14929_/A sky130_fd_sc_hd__and2_1
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14858_ hold17/A _16303_/Q hold19/A _14818_/X vssd1 vssd1 vccd1 vccd1 _16287_/D sky130_fd_sc_hd__o31a_1
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13809_ _13809_/A _13809_/B vssd1 vssd1 vccd1 vccd1 _13812_/C sky130_fd_sc_hd__nor2_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14789_ _14988_/A vssd1 vssd1 vccd1 vccd1 _14789_/X sky130_fd_sc_hd__buf_2
XFILLER_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09000_ _09000_/A vssd1 vssd1 vccd1 vccd1 _15302_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09902_ _09902_/A vssd1 vssd1 vccd1 vccd1 _15442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09833_ _15431_/Q vssd1 vssd1 vccd1 vccd1 _09847_/C sky130_fd_sc_hd__inv_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09764_ _09997_/A _09764_/B _09764_/C vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__or3_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08715_ _15260_/Q _08775_/B _08715_/C vssd1 vssd1 vccd1 vccd1 _08724_/B sky130_fd_sc_hd__and3_1
X_09695_ _15410_/Q _09813_/B _09700_/C vssd1 vssd1 vccd1 vccd1 _09695_/Y sky130_fd_sc_hd__nand3_1
XFILLER_54_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08646_ _08643_/X _08644_/Y _08645_/Y _08639_/C vssd1 vssd1 vccd1 vccd1 _08648_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ hold36/X _10957_/C _08582_/C vssd1 vssd1 vccd1 vccd1 _08577_/Y sky130_fd_sc_hd__nand3_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ _10484_/C vssd1 vssd1 vccd1 vccd1 _10492_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09129_ _09129_/A _09129_/B vssd1 vssd1 vccd1 vccd1 _09133_/C sky130_fd_sc_hd__nor2_1
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12140_ _15793_/Q _12178_/C _11912_/X vssd1 vssd1 vccd1 vccd1 _12142_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _12639_/A vssd1 vssd1 vccd1 vccd1 _12299_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _15618_/Q _11027_/C _10848_/X vssd1 vssd1 vccd1 vccd1 _11022_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15830_ _07603_/A _15830_/D vssd1 vssd1 vccd1 vccd1 _15830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15761_ _15763_/CLK _15761_/D vssd1 vssd1 vccd1 vccd1 _15761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12973_ _12973_/A _12973_/B vssd1 vssd1 vccd1 vccd1 _12977_/C sky130_fd_sc_hd__nor2_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14712_ _16258_/Q _14833_/B _14717_/C vssd1 vssd1 vccd1 vccd1 _14721_/A sky130_fd_sc_hd__and3_1
XFILLER_18_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11924_ _15759_/Q _11931_/C _11805_/X vssd1 vssd1 vccd1 vccd1 _11924_/Y sky130_fd_sc_hd__a21oi_1
X_15692_ _15692_/CLK _15692_/D vssd1 vssd1 vccd1 vccd1 _15692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14643_ _14643_/A _14643_/B vssd1 vssd1 vccd1 vccd1 _14644_/B sky130_fd_sc_hd__nor2_1
X_11855_ _11949_/A _11855_/B _11860_/A vssd1 vssd1 vccd1 vccd1 _15747_/D sky130_fd_sc_hd__nor3_1
XFILLER_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10806_ _10863_/A _10806_/B _10806_/C vssd1 vssd1 vccd1 vccd1 _10808_/B sky130_fd_sc_hd__or3_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14574_ _14408_/X _14572_/B _14573_/Y vssd1 vssd1 vccd1 vccd1 _16221_/D sky130_fd_sc_hd__o21a_1
X_11786_ _11824_/A _11786_/B _11786_/C vssd1 vssd1 vccd1 vccd1 _11787_/A sky130_fd_sc_hd__and3_1
X_16313_ _16327_/CLK _16313_/D vssd1 vssd1 vccd1 vccd1 _16313_/Q sky130_fd_sc_hd__dfxtp_1
X_13525_ _16021_/Q _13628_/B _13533_/C vssd1 vssd1 vccd1 vccd1 _13529_/B sky130_fd_sc_hd__nand3_1
X_10737_ _15572_/Q _11023_/B _10741_/C vssd1 vssd1 vccd1 vccd1 _10737_/Y sky130_fd_sc_hd__nand3_1
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16244_ _16264_/CLK _16244_/D vssd1 vssd1 vccd1 vccd1 _16244_/Q sky130_fd_sc_hd__dfxtp_2
X_13456_ _13456_/A _13456_/B vssd1 vssd1 vccd1 vccd1 _13460_/C sky130_fd_sc_hd__nor2_1
XFILLER_139_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10668_ _10676_/A _10668_/B _10668_/C vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__and3_1
X_12407_ _12414_/B _12407_/B vssd1 vssd1 vccd1 vccd1 _12410_/A sky130_fd_sc_hd__or2_1
XFILLER_126_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16175_ _16192_/CLK _16175_/D vssd1 vssd1 vccd1 vccd1 _16175_/Q sky130_fd_sc_hd__dfxtp_1
X_10599_ _10593_/B _10594_/C _10596_/X _10597_/Y vssd1 vssd1 vccd1 vccd1 _10600_/C
+ sky130_fd_sc_hd__a211o_1
X_13387_ _15996_/Q _13589_/B _13394_/C vssd1 vssd1 vccd1 vccd1 _13387_/X sky130_fd_sc_hd__and3_1
XFILLER_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15126_ _16341_/Q vssd1 vssd1 vccd1 vccd1 _15131_/C sky130_fd_sc_hd__inv_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12338_ _12338_/A vssd1 vssd1 vccd1 vccd1 _15823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15057_ _15061_/C vssd1 vssd1 vccd1 vccd1 _15072_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12269_ _15814_/Q _12270_/C _12100_/X vssd1 vssd1 vccd1 vccd1 _12269_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14008_ _14002_/Y _14006_/X _14007_/Y vssd1 vssd1 vccd1 vccd1 _16103_/D sky130_fd_sc_hd__o21a_1
XFILLER_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15959_ _15970_/CLK _15959_/D vssd1 vssd1 vccd1 vccd1 _15959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08500_ _15230_/Q _11128_/A _08505_/C vssd1 vssd1 vccd1 vccd1 _08500_/X sky130_fd_sc_hd__and3_1
X_09480_ _15385_/Q _15384_/Q _15383_/Q _09194_/X vssd1 vssd1 vccd1 vccd1 _15377_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_64_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08431_ _08428_/Y _08430_/Y _08168_/X vssd1 vssd1 vccd1 vccd1 _08431_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08362_ _08362_/A _08362_/B vssd1 vssd1 vccd1 vccd1 _08363_/B sky130_fd_sc_hd__xnor2_2
XFILLER_32_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08293_ _08293_/A _08293_/B vssd1 vssd1 vccd1 vccd1 _08296_/A sky130_fd_sc_hd__nand2_2
XFILLER_149_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09816_ _09930_/A _09816_/B _09820_/B vssd1 vssd1 vccd1 vccd1 _15428_/D sky130_fd_sc_hd__nor3_1
XFILLER_59_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09747_ _09747_/A vssd1 vssd1 vccd1 vccd1 _15418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _15409_/Q _09680_/C _09506_/X vssd1 vssd1 vccd1 vccd1 _09678_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08648_/A _08629_/B _08629_/C vssd1 vssd1 vccd1 vccd1 _08630_/A sky130_fd_sc_hd__and3_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11640_ _11640_/A vssd1 vssd1 vccd1 vccd1 _15713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ _15704_/Q _11576_/C _11512_/X vssd1 vssd1 vccd1 vccd1 _11573_/C sky130_fd_sc_hd__a21o_1
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13310_ _13153_/X _13307_/C _13309_/Y vssd1 vssd1 vccd1 vccd1 _15980_/D sky130_fd_sc_hd__a21oi_1
X_10522_ _10559_/A _10522_/B _10522_/C vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__and3_1
X_14290_ _14304_/A _14290_/B _14295_/A vssd1 vssd1 vccd1 vccd1 _16162_/D sky130_fd_sc_hd__nor3_1
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10453_ _15529_/Q _10512_/B _10453_/C vssd1 vssd1 vccd1 vccd1 _10463_/B sky130_fd_sc_hd__and3_1
XFILLER_108_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13241_ _15970_/Q _13246_/C _14605_/B vssd1 vssd1 vccd1 vccd1 _13241_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10384_ _10381_/X _10382_/Y _10383_/Y _10378_/C vssd1 vssd1 vccd1 vccd1 _10386_/B
+ sky130_fd_sc_hd__o211ai_1
X_13172_ _15959_/Q _14298_/A _13172_/C vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__and3_1
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ _12130_/B _12123_/B vssd1 vssd1 vccd1 vccd1 _12126_/A sky130_fd_sc_hd__or2_1
X_12054_ _12054_/A vssd1 vssd1 vccd1 vccd1 _15778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11005_ _11582_/A vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_77_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15813_ _07603_/A _15813_/D vssd1 vssd1 vccd1 vccd1 _15813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15744_ _15763_/CLK _15744_/D vssd1 vssd1 vccd1 vccd1 _15744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12956_ _15922_/Q _13066_/B _12962_/C vssd1 vssd1 vccd1 vccd1 _12956_/Y sky130_fd_sc_hd__nand3_1
XFILLER_18_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11907_ _15755_/Q vssd1 vssd1 vccd1 vccd1 _11923_/C sky130_fd_sc_hd__inv_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _15763_/CLK _15675_/D vssd1 vssd1 vccd1 vccd1 _15675_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12887_ _15912_/Q _12996_/B _12887_/C vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__and3_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14626_ _14626_/A _14626_/B _14630_/A vssd1 vssd1 vccd1 vccd1 _16234_/D sky130_fd_sc_hd__nor3_1
X_11838_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12068_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14551_/B _14552_/C _14561_/A _14555_/Y vssd1 vssd1 vccd1 vccd1 _14561_/B
+ sky130_fd_sc_hd__a211oi_1
X_11769_ _15734_/Q _11887_/B _11774_/C vssd1 vssd1 vccd1 vccd1 _11769_/Y sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_40_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16169_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _14879_/A vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14488_ _14486_/X _14488_/B vssd1 vssd1 vccd1 vccd1 _14488_/X sky130_fd_sc_hd__and2b_1
X_16227_ _16241_/CLK _16227_/D vssd1 vssd1 vccd1 vccd1 _16227_/Q sky130_fd_sc_hd__dfxtp_2
X_13439_ _16004_/Q _13543_/B _13445_/C vssd1 vssd1 vccd1 vccd1 _13439_/Y sky130_fd_sc_hd__nand3_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16158_ _16169_/CLK _16158_/D vssd1 vssd1 vccd1 vccd1 _16158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15109_ _15109_/A _15109_/B vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__or2_1
X_08980_ _10134_/A vssd1 vssd1 vccd1 vccd1 _09211_/B sky130_fd_sc_hd__clkbuf_4
X_16089_ _16119_/CLK _16089_/D vssd1 vssd1 vccd1 vccd1 _16089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07931_ _15342_/Q _07932_/B vssd1 vssd1 vccd1 vccd1 _07933_/A sky130_fd_sc_hd__or2_1
XFILLER_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07862_ _15818_/Q vssd1 vssd1 vccd1 vccd1 _12304_/A sky130_fd_sc_hd__inv_2
XFILLER_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09601_ _09601_/A vssd1 vssd1 vccd1 vccd1 _09615_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07793_ _16224_/Q vssd1 vssd1 vccd1 vccd1 _08065_/A sky130_fd_sc_hd__inv_2
XFILLER_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09532_ _10110_/A vssd1 vssd1 vccd1 vccd1 _09760_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09463_ _09470_/A _09461_/Y _09462_/Y _09458_/C vssd1 vssd1 vccd1 vccd1 _09465_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08414_ _08414_/A _08414_/B vssd1 vssd1 vccd1 vccd1 _08414_/X sky130_fd_sc_hd__or2_1
X_09394_ _09401_/A _09394_/B _09394_/C vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__and3_1
X_08345_ _08384_/A _08384_/C vssd1 vssd1 vccd1 vccd1 _08346_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_31_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15935_/CLK sky130_fd_sc_hd__clkbuf_16
X_08276_ _07946_/C _08166_/Y _08275_/X vssd1 vssd1 vccd1 vccd1 _08276_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12810_ _12919_/A _12813_/C vssd1 vssd1 vccd1 vccd1 _12810_/X sky130_fd_sc_hd__or2_1
XFILLER_90_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13790_ _13790_/A vssd1 vssd1 vccd1 vccd1 _16065_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12741_/A vssd1 vssd1 vccd1 vccd1 _15886_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _15483_/CLK _15460_/D vssd1 vssd1 vccd1 vccd1 _15460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12670_/Y _12665_/C _12667_/X _12669_/Y vssd1 vssd1 vccd1 vccd1 _12673_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14411_ _14533_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14411_/Y sky130_fd_sc_hd__nor2_1
X_11623_ _11655_/C vssd1 vssd1 vccd1 vccd1 _11662_/C sky130_fd_sc_hd__clkbuf_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _15484_/CLK _15391_/D vssd1 vssd1 vccd1 vccd1 _15391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _16075_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14342_ _14342_/A _14342_/B _14342_/C vssd1 vssd1 vccd1 vccd1 _14343_/C sky130_fd_sc_hd__nand3_1
X_11554_ _11552_/A _11552_/B _11553_/X vssd1 vssd1 vccd1 vccd1 _15699_/D sky130_fd_sc_hd__a21oi_1
XFILLER_11_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10505_ _11422_/A vssd1 vssd1 vccd1 vccd1 _10734_/B sky130_fd_sc_hd__clkbuf_2
X_14273_ _14268_/Y _14272_/X _14196_/X vssd1 vssd1 vccd1 vccd1 _14273_/Y sky130_fd_sc_hd__a21oi_1
X_11485_ input7/X vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__buf_2
XFILLER_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16012_ _16022_/CLK _16012_/D vssd1 vssd1 vccd1 vccd1 _16012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13224_ _13224_/A vssd1 vssd1 vccd1 vccd1 _15965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ _10434_/Y _10430_/C _10432_/X _10433_/Y vssd1 vssd1 vccd1 vccd1 _10437_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13155_ _13154_/X _13149_/C _08335_/X vssd1 vssd1 vccd1 vccd1 _13155_/Y sky130_fd_sc_hd__o21ai_1
X_10367_ _10360_/B _10361_/C _10363_/X _10365_/Y vssd1 vssd1 vccd1 vccd1 _10368_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _12106_/A vssd1 vssd1 vccd1 vccd1 _15786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10298_ _15506_/Q _10298_/B _10304_/C vssd1 vssd1 vccd1 vccd1 _10301_/B sky130_fd_sc_hd__nand3_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13086_ _13151_/A _13086_/B _13086_/C vssd1 vssd1 vccd1 vccd1 _13088_/B sky130_fd_sc_hd__or3_1
XFILLER_78_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_89_clk _15584_/CLK vssd1 vssd1 vccd1 vccd1 _15239_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12037_ _12053_/A _12037_/B _12037_/C vssd1 vssd1 vccd1 vccd1 _12038_/A sky130_fd_sc_hd__and3_1
XFILLER_120_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13988_ _14541_/A vssd1 vssd1 vccd1 vccd1 _14434_/A sky130_fd_sc_hd__buf_4
X_15727_ _15763_/CLK _15727_/D vssd1 vssd1 vccd1 vccd1 _15727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12939_ _12959_/A _12939_/B _12939_/C vssd1 vssd1 vccd1 vccd1 _12940_/A sky130_fd_sc_hd__and3_1
XFILLER_34_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15658_ _15763_/CLK _15658_/D vssd1 vssd1 vccd1 vccd1 _15658_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14609_ _14604_/Y _14607_/X _14608_/Y vssd1 vssd1 vccd1 vccd1 _16229_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15589_ _15194_/Q _15589_/D vssd1 vssd1 vccd1 vccd1 _15589_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_13_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _16011_/CLK sky130_fd_sc_hd__clkbuf_16
X_08130_ _08243_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _08131_/B sky130_fd_sc_hd__xnor2_2
XFILLER_119_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08061_ _08062_/A _08062_/B vssd1 vssd1 vccd1 vccd1 _08211_/B sky130_fd_sc_hd__nor2_1
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08963_ _08999_/A _08963_/B _08963_/C vssd1 vssd1 vccd1 vccd1 _08964_/A sky130_fd_sc_hd__and3_1
XFILLER_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07914_ hold28/A _16305_/Q vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08894_ _08892_/A _08892_/B _08893_/X vssd1 vssd1 vccd1 vccd1 _15286_/D sky130_fd_sc_hd__a21oi_1
XFILLER_111_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07845_ _15854_/Q _08022_/B vssd1 vssd1 vccd1 vccd1 _07846_/B sky130_fd_sc_hd__xnor2_4
XFILLER_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07776_ _07777_/A _07778_/B vssd1 vssd1 vccd1 vccd1 _07779_/A sky130_fd_sc_hd__or2_1
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09515_ _15383_/Q _09522_/C _09453_/X vssd1 vssd1 vccd1 vccd1 _09515_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _15372_/Q _09623_/B _09446_/C vssd1 vssd1 vccd1 vccd1 _09446_/Y sky130_fd_sc_hd__nand3_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09377_ _09377_/A _09377_/B _09377_/C vssd1 vssd1 vccd1 vccd1 _09378_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08328_ _08365_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__or2_1
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08259_ _08259_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__xnor2_4
XFILLER_119_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11270_ _11309_/A _11270_/B _11270_/C vssd1 vssd1 vccd1 vccd1 _11271_/A sky130_fd_sc_hd__and3_1
X_10221_ _15493_/Q _10220_/C _10044_/X vssd1 vssd1 vccd1 vccd1 _10222_/B sky130_fd_sc_hd__a21oi_1
XFILLER_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10152_ _10150_/Y _10146_/C _10148_/X _10149_/Y vssd1 vssd1 vccd1 vccd1 _10153_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_121_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10083_ _10663_/A vssd1 vssd1 vccd1 vccd1 _10083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14960_ _14955_/A _14958_/B _14845_/X vssd1 vssd1 vccd1 vccd1 _14967_/C sky130_fd_sc_hd__o21a_1
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _15189_/A vssd1 vssd1 vccd1 vccd1 _14408_/A sky130_fd_sc_hd__buf_2
XFILLER_75_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14891_ _15051_/A _15010_/B _14891_/C vssd1 vssd1 vccd1 vccd1 _14895_/A sky130_fd_sc_hd__and3_1
XFILLER_114_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13842_ _13838_/X _13839_/Y _13841_/Y _13836_/C vssd1 vssd1 vccd1 vccd1 _13844_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13773_ _13777_/C vssd1 vssd1 vccd1 vccd1 _13785_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10985_ _15611_/Q vssd1 vssd1 vccd1 vccd1 _10999_/C sky130_fd_sc_hd__inv_2
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15512_ _15512_/CLK _15512_/D vssd1 vssd1 vccd1 vccd1 _15512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12724_ _12740_/A _12724_/B _12724_/C vssd1 vssd1 vccd1 vccd1 _12725_/A sky130_fd_sc_hd__and3_1
XFILLER_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15443_ _15483_/CLK _15443_/D vssd1 vssd1 vccd1 vccd1 _15443_/Q sky130_fd_sc_hd__dfxtp_1
X_12655_ _15875_/Q _12660_/C _12654_/X vssd1 vssd1 vccd1 vccd1 _12657_/C sky130_fd_sc_hd__a21o_1
X_11606_ _15709_/Q _11605_/C _11488_/X vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__a21oi_1
X_15374_ _15484_/CLK _15374_/D vssd1 vssd1 vccd1 vccd1 _15374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12586_ _12586_/A vssd1 vssd1 vccd1 vccd1 _15862_/D sky130_fd_sc_hd__clkbuf_1
X_14325_ _14325_/A vssd1 vssd1 vccd1 vccd1 _14325_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11537_ _11535_/Y _11531_/C _11533_/X _11534_/Y vssd1 vssd1 vccd1 vccd1 _11538_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14256_ _16158_/Q _14256_/B _14256_/C vssd1 vssd1 vccd1 vccd1 _14264_/A sky130_fd_sc_hd__and3_1
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11468_ _11466_/Y _11461_/C _11463_/X _11464_/Y vssd1 vssd1 vccd1 vccd1 _11469_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_109_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13207_ _13154_/X _13204_/C _13206_/X vssd1 vssd1 vccd1 vccd1 _13207_/Y sky130_fd_sc_hd__o21ai_1
X_10419_ _15524_/Q _10426_/C _10357_/X vssd1 vssd1 vccd1 vccd1 _10421_/C sky130_fd_sc_hd__a21o_1
XFILLER_99_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14187_ _14185_/X _14187_/B vssd1 vssd1 vccd1 vccd1 _14187_/X sky130_fd_sc_hd__and2b_1
X_11399_ _11420_/A _11399_/B _11399_/C vssd1 vssd1 vccd1 vccd1 _11400_/A sky130_fd_sc_hd__and3_1
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _15953_/Q _13349_/B _13138_/C vssd1 vssd1 vccd1 vccd1 _13146_/B sky130_fd_sc_hd__and3_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _13069_/A _13069_/B _13069_/C vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__and3_1
XFILLER_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_clk _15665_/CLK vssd1 vssd1 vccd1 vccd1 _15620_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07630_ _13045_/B vssd1 vssd1 vccd1 vccd1 _07634_/A sky130_fd_sc_hd__buf_6
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09300_ _09300_/A _09300_/B vssd1 vssd1 vccd1 vccd1 _09301_/B sky130_fd_sc_hd__nor2_1
XFILLER_62_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09231_ _09228_/X _09229_/Y _09230_/Y _09225_/C vssd1 vssd1 vccd1 vccd1 _09233_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09162_ _09160_/Y _09156_/C _09158_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _09163_/C
+ sky130_fd_sc_hd__a211o_1
X_08113_ _15413_/Q _08113_/B vssd1 vssd1 vccd1 vccd1 _08113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09093_ _09093_/A _09093_/B _09093_/C vssd1 vssd1 vccd1 vccd1 _09094_/C sky130_fd_sc_hd__nand3_1
X_08044_ _08044_/A _07823_/B vssd1 vssd1 vccd1 vccd1 _08044_/X sky130_fd_sc_hd__or2b_1
XFILLER_115_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09995_ _09993_/A _09993_/B _09994_/X vssd1 vssd1 vccd1 vccd1 _15456_/D sky130_fd_sc_hd__a21oi_1
XFILLER_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08946_ _15295_/Q _08951_/C _08824_/X vssd1 vssd1 vccd1 vccd1 _08946_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08877_ _08875_/Y _08870_/C _08872_/X _08874_/Y vssd1 vssd1 vccd1 vccd1 _08878_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07828_ _07828_/A _07828_/B vssd1 vssd1 vccd1 vccd1 _08148_/B sky130_fd_sc_hd__xor2_4
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07759_ _15692_/Q vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__clkinv_4
X_10770_ _15579_/Q _10999_/B _10770_/C vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__and3_1
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09429_ _10007_/A vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12440_ _12726_/A vssd1 vssd1 vccd1 vccd1 _12667_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_60_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12371_ _15830_/Q _12376_/C _12370_/X vssd1 vssd1 vccd1 vccd1 _12373_/C sky130_fd_sc_hd__a21o_1
X_14110_ _13666_/A _14108_/C _13720_/X vssd1 vssd1 vccd1 vccd1 _14110_/Y sky130_fd_sc_hd__o21ai_1
X_11322_ _11493_/A _11326_/C vssd1 vssd1 vccd1 vccd1 _11322_/X sky130_fd_sc_hd__or2_1
X_15090_ _15013_/X _15088_/A _15089_/Y vssd1 vssd1 vccd1 vccd1 _16340_/D sky130_fd_sc_hd__o21a_1
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14041_ _14041_/A _14041_/B vssd1 vssd1 vccd1 vccd1 _14041_/X sky130_fd_sc_hd__or2_1
X_11253_ _15654_/Q _11367_/B _11253_/C vssd1 vssd1 vccd1 vccd1 _11262_/A sky130_fd_sc_hd__and3_1
XFILLER_134_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10204_ _15491_/Q _10317_/B _10214_/C vssd1 vssd1 vccd1 vccd1 _10204_/X sky130_fd_sc_hd__and3_1
X_11184_ _12048_/A vssd1 vssd1 vccd1 vccd1 _11184_/X sky130_fd_sc_hd__buf_2
XFILLER_122_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10135_ _15480_/Q _10363_/B _10135_/C vssd1 vssd1 vccd1 vccd1 _10135_/X sky130_fd_sc_hd__and3_1
XFILLER_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15992_ _15994_/CLK _15992_/D vssd1 vssd1 vccd1 vccd1 _15992_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10066_ _15470_/Q _10298_/B _10074_/C vssd1 vssd1 vccd1 vccd1 _10071_/B sky130_fd_sc_hd__nand3_1
X_14943_ _16311_/Q _14941_/C _14942_/X vssd1 vssd1 vccd1 vccd1 _14945_/C sky130_fd_sc_hd__a21o_1
XFILLER_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14874_ _14915_/A _14874_/B _14878_/B vssd1 vssd1 vccd1 vccd1 _16290_/D sky130_fd_sc_hd__nor3_1
XFILLER_36_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13825_ _13852_/A _13825_/B _13829_/A vssd1 vssd1 vccd1 vccd1 _16072_/D sky130_fd_sc_hd__nor3_1
XFILLER_90_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13756_ _13754_/Y _13749_/C _13761_/A _13753_/Y vssd1 vssd1 vccd1 vccd1 _13761_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10968_ _11085_/A _10968_/B _10973_/B vssd1 vssd1 vccd1 vccd1 _15608_/D sky130_fd_sc_hd__nor3_1
XFILLER_71_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12707_ _12720_/C vssd1 vssd1 vccd1 vccd1 _12729_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13687_ _16049_/Q _13686_/C _13534_/X vssd1 vssd1 vccd1 vccd1 _13687_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10899_ _15598_/Q _11073_/B _10904_/C vssd1 vssd1 vccd1 vccd1 _10899_/Y sky130_fd_sc_hd__nand3_1
X_15426_ _15483_/CLK _15426_/D vssd1 vssd1 vccd1 vccd1 _15426_/Q sky130_fd_sc_hd__dfxtp_1
X_12638_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12680_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15357_ _15359_/CLK _15357_/D vssd1 vssd1 vccd1 vccd1 _15357_/Q sky130_fd_sc_hd__dfxtp_1
X_12569_ _12569_/A vssd1 vssd1 vccd1 vccd1 _12569_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14308_ _14308_/A _14308_/B vssd1 vssd1 vccd1 vccd1 _14308_/X sky130_fd_sc_hd__or2_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15288_ _16344_/CLK _15288_/D vssd1 vssd1 vccd1 vccd1 _15288_/Q sky130_fd_sc_hd__dfxtp_1
X_14239_ _14058_/X _14235_/B _14059_/X vssd1 vssd1 vccd1 vccd1 _14242_/A sky130_fd_sc_hd__a21oi_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08821_/A _08800_/B _08800_/C vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__and3_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09781_/B _09781_/C _09781_/A vssd1 vssd1 vccd1 vccd1 _09782_/B sky130_fd_sc_hd__a21o_1
XFILLER_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08745_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08662_ _14541_/A vssd1 vssd1 vccd1 vccd1 _08893_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07613_ _15030_/A vssd1 vssd1 vccd1 vccd1 _08421_/A sky130_fd_sc_hd__clkbuf_4
X_08593_ _08593_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _08594_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09214_ _09211_/X _09213_/Y _09208_/B _09209_/C vssd1 vssd1 vccd1 vccd1 _09216_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_139_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ _09202_/A _09145_/B _09149_/A vssd1 vssd1 vccd1 vccd1 _15325_/D sky130_fd_sc_hd__nor3_1
X_09076_ _09075_/B _09075_/C _09019_/X vssd1 vssd1 vccd1 vccd1 _09077_/C sky130_fd_sc_hd__o21ai_1
XFILLER_108_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08027_ _14380_/C _08027_/B vssd1 vssd1 vccd1 vccd1 _08033_/A sky130_fd_sc_hd__or2_1
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09978_ _09978_/A vssd1 vssd1 vccd1 vccd1 _15454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08929_ _13057_/B vssd1 vssd1 vccd1 vccd1 _08929_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11940_ _11938_/Y _11934_/C _11936_/X _11937_/Y vssd1 vssd1 vccd1 vccd1 _11941_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11871_ _15751_/Q _11872_/C _11812_/X vssd1 vssd1 vccd1 vccd1 _11871_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13610_ _13713_/A _13613_/C vssd1 vssd1 vccd1 vccd1 _13610_/X sky130_fd_sc_hd__or2_1
X_10822_ _10822_/A _10822_/B _10822_/C vssd1 vssd1 vccd1 vccd1 _10823_/C sky130_fd_sc_hd__nand3_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14590_ _14590_/A _14590_/B _14590_/C vssd1 vssd1 vccd1 vccd1 _14591_/C sky130_fd_sc_hd__nand3_1
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13541_ _16023_/Q _13589_/B _13548_/C vssd1 vssd1 vccd1 vccd1 _13541_/X sky130_fd_sc_hd__and3_1
X_10753_ _10789_/A _10753_/B _10753_/C vssd1 vssd1 vccd1 vccd1 _10754_/A sky130_fd_sc_hd__and3_1
XFILLER_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16260_ _16317_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 _16260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13472_ _13498_/C vssd1 vssd1 vccd1 vccd1 _13504_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10684_ _10797_/A _10684_/B _10688_/B vssd1 vssd1 vccd1 vccd1 _15563_/D sky130_fd_sc_hd__nor3_1
XFILLER_139_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15211_ _16353_/CLK _15211_/D vssd1 vssd1 vccd1 vccd1 _15211_/Q sky130_fd_sc_hd__dfxtp_1
X_12423_ _12456_/C vssd1 vssd1 vccd1 vccd1 _12462_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16191_ _16247_/CLK _16191_/D vssd1 vssd1 vccd1 vccd1 _16191_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15142_ _16358_/Q _15142_/B _15142_/C vssd1 vssd1 vccd1 vccd1 _15144_/A sky130_fd_sc_hd__and3_1
X_12354_ _12413_/A vssd1 vssd1 vccd1 vccd1 _12396_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ _15662_/Q _11311_/C _11184_/X vssd1 vssd1 vccd1 vccd1 _11305_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15073_ hold15/X _15072_/C _14917_/X vssd1 vssd1 vccd1 vccd1 _15074_/B sky130_fd_sc_hd__a21oi_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12285_ _12569_/A vssd1 vssd1 vccd1 vccd1 _12285_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ _14291_/A vssd1 vssd1 vccd1 vccd1 _14249_/B sky130_fd_sc_hd__buf_2
X_11236_ _15652_/Q _11236_/B _11239_/C vssd1 vssd1 vccd1 vccd1 _11236_/X sky130_fd_sc_hd__and3_1
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11167_ _11189_/A _11167_/B _11167_/C vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__and3_1
XFILLER_121_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10118_ _10118_/A vssd1 vssd1 vccd1 vccd1 _15475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11098_ _15637_/Q _15636_/Q _15635_/Q _10983_/X vssd1 vssd1 vccd1 vccd1 _15629_/D
+ sky130_fd_sc_hd__o31a_1
X_15975_ _15984_/CLK _15975_/D vssd1 vssd1 vccd1 vccd1 _15975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10049_ _10049_/A _10053_/C vssd1 vssd1 vccd1 vccd1 _10049_/X sky130_fd_sc_hd__or2_1
X_14926_ _14802_/X _14919_/A _14922_/B _14925_/Y vssd1 vssd1 vccd1 vccd1 _16301_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_75_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14857_ _14814_/X _14855_/A _14856_/Y vssd1 vssd1 vccd1 vccd1 _16286_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13808_ _13808_/A _13808_/B vssd1 vssd1 vccd1 vccd1 _13809_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14788_ hold14/A _14833_/B _14795_/C vssd1 vssd1 vccd1 vccd1 _14798_/A sky130_fd_sc_hd__and3_1
XFILLER_51_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13739_ _16058_/Q _13738_/C _13534_/X vssd1 vssd1 vccd1 vccd1 _13739_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ _15483_/CLK _15409_/D vssd1 vssd1 vccd1 vccd1 _15409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ _09922_/A _09901_/B _09901_/C vssd1 vssd1 vccd1 vccd1 _09902_/A sky130_fd_sc_hd__and3_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _15439_/Q _15438_/Q _15437_/Q _09831_/X vssd1 vssd1 vccd1 vccd1 _15431_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _10341_/A vssd1 vssd1 vccd1 vccd1 _09997_/A sky130_fd_sc_hd__clkbuf_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08714_ _08774_/A _08714_/B _08718_/B vssd1 vssd1 vccd1 vccd1 _15258_/D sky130_fd_sc_hd__nor3_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09694_ _15411_/Q _09700_/C _09693_/X vssd1 vssd1 vccd1 vccd1 _09694_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _15248_/Q _10957_/C _08651_/C vssd1 vssd1 vccd1 vccd1 _08645_/Y sky130_fd_sc_hd__nand3_1
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08576_ _15240_/Q _08582_/C _08575_/X vssd1 vssd1 vccd1 vccd1 _08576_/Y sky130_fd_sc_hd__a21oi_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09128_ _09128_/A _09128_/B vssd1 vssd1 vccd1 vccd1 _09129_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09059_ _09059_/A vssd1 vssd1 vccd1 vccd1 _15311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12070_ _12129_/A vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11021_ _15618_/Q _11078_/B _11021_/C vssd1 vssd1 vccd1 vccd1 _11030_/A sky130_fd_sc_hd__and3_1
XFILLER_103_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15760_ _15794_/CLK _15760_/D vssd1 vssd1 vccd1 vccd1 _15760_/Q sky130_fd_sc_hd__dfxtp_1
X_12972_ _12972_/A vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11923_ _15759_/Q _12150_/B _11923_/C vssd1 vssd1 vccd1 vccd1 _11923_/X sky130_fd_sc_hd__and3_1
X_14711_ _14711_/A vssd1 vssd1 vccd1 vccd1 _16253_/D sky130_fd_sc_hd__clkbuf_1
X_15691_ _15763_/CLK _15691_/D vssd1 vssd1 vccd1 vccd1 _15691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14642_ _14642_/A _14642_/B vssd1 vssd1 vccd1 vccd1 _14643_/B sky130_fd_sc_hd__nor2_1
X_11854_ _15748_/Q _12025_/B _11863_/C vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__and3_1
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10805_ _10978_/A vssd1 vssd1 vccd1 vccd1 _10845_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14573_ _14612_/A _14573_/B vssd1 vssd1 vccd1 vccd1 _14573_/Y sky130_fd_sc_hd__nor2_1
X_11785_ _11784_/B _11784_/C _11615_/X vssd1 vssd1 vccd1 vccd1 _11786_/C sky130_fd_sc_hd__o21ai_1
XFILLER_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16312_ _16312_/CLK _16312_/D vssd1 vssd1 vccd1 vccd1 _16312_/Q sky130_fd_sc_hd__dfxtp_1
X_13524_ _13604_/A _13524_/B _13529_/A vssd1 vssd1 vccd1 vccd1 _16018_/D sky130_fd_sc_hd__nor3_1
X_10736_ _10736_/A vssd1 vssd1 vccd1 vccd1 _11023_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16243_ _16247_/CLK _16243_/D vssd1 vssd1 vccd1 vccd1 _16243_/Q sky130_fd_sc_hd__dfxtp_2
X_13455_ _13455_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13456_/B sky130_fd_sc_hd__nor2_1
X_10667_ _10665_/Y _10659_/C _10662_/X _10664_/Y vssd1 vssd1 vccd1 vccd1 _10668_/C
+ sky130_fd_sc_hd__a211o_1
X_12406_ _15835_/Q _12405_/C _12347_/X vssd1 vssd1 vccd1 vccd1 _12407_/B sky130_fd_sc_hd__a21oi_1
X_16174_ _16187_/CLK _16174_/D vssd1 vssd1 vccd1 vccd1 _16174_/Q sky130_fd_sc_hd__dfxtp_1
X_13386_ _13640_/A vssd1 vssd1 vccd1 vccd1 _13589_/B sky130_fd_sc_hd__clkbuf_4
X_10598_ _10596_/X _10597_/Y _10593_/B _10594_/C vssd1 vssd1 vccd1 vccd1 _10600_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_126_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15125_ _16367_/Q _16366_/Q _16365_/Q _15017_/X vssd1 vssd1 vccd1 vccd1 _16350_/D
+ sky130_fd_sc_hd__o31a_1
X_12337_ _12337_/A _12337_/B _12337_/C vssd1 vssd1 vccd1 vccd1 _12338_/A sky130_fd_sc_hd__and3_1
XFILLER_114_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15056_ _16349_/Q _16348_/Q _16347_/Q _15017_/X vssd1 vssd1 vccd1 vccd1 _16332_/D
+ sky130_fd_sc_hd__o31a_1
X_12268_ _15814_/Q _12383_/B _12270_/C vssd1 vssd1 vccd1 vccd1 _12268_/X sky130_fd_sc_hd__and3_1
XFILLER_142_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14007_ _14002_/Y _14006_/X _13922_/X vssd1 vssd1 vccd1 vccd1 _14007_/Y sky130_fd_sc_hd__a21oi_1
X_11219_ _15649_/Q _11449_/B _11228_/C vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__and3_1
X_12199_ _15802_/Q _12309_/B _12208_/C vssd1 vssd1 vccd1 vccd1 _12204_/A sky130_fd_sc_hd__and3_1
XFILLER_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15958_ _15970_/CLK _15958_/D vssd1 vssd1 vccd1 vccd1 _15958_/Q sky130_fd_sc_hd__dfxtp_1
X_14909_ _14946_/A _14909_/B _14909_/C vssd1 vssd1 vccd1 vccd1 _14910_/A sky130_fd_sc_hd__and3_1
X_15889_ _07603_/A _15889_/D vssd1 vssd1 vccd1 vccd1 _15889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08430_ _08421_/C _08424_/Y _08429_/X vssd1 vssd1 vccd1 vccd1 _08430_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08361_ _08381_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _08362_/B sky130_fd_sc_hd__xor2_2
XFILLER_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08292_ _08292_/A _08194_/A vssd1 vssd1 vccd1 vccd1 _08293_/B sky130_fd_sc_hd__or2b_1
XFILLER_20_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09815_ _09813_/Y _09807_/C _09820_/A _09812_/Y vssd1 vssd1 vccd1 vccd1 _09820_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09746_ _09746_/A _09746_/B _09746_/C vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__and3_1
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _15409_/Q _09733_/B _09680_/C vssd1 vssd1 vccd1 vccd1 _09677_/X sky130_fd_sc_hd__and3_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _08619_/B _08620_/C _08622_/X _08626_/Y vssd1 vssd1 vccd1 vccd1 _08629_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08559_/A vssd1 vssd1 vccd1 vccd1 _15236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11570_ _15704_/Q _11797_/B _11576_/C vssd1 vssd1 vccd1 vccd1 _11573_/B sky130_fd_sc_hd__nand3_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10521_ _10520_/B _10520_/C _10464_/X vssd1 vssd1 vccd1 vccd1 _10522_/C sky130_fd_sc_hd__o21ai_1
XFILLER_149_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _15970_/Q _13394_/B _13240_/C vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__and3_1
X_10452_ _10511_/A _10452_/B _10456_/B vssd1 vssd1 vccd1 vccd1 _15527_/D sky130_fd_sc_hd__nor3_1
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ _13171_/A vssd1 vssd1 vccd1 vccd1 _15956_/D sky130_fd_sc_hd__clkbuf_1
X_10383_ _15517_/Q _10441_/B _10389_/C vssd1 vssd1 vccd1 vccd1 _10383_/Y sky130_fd_sc_hd__nand3_1
XFILLER_123_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12122_ _15790_/Q _12121_/C _12063_/X vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__a21oi_1
XFILLER_124_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12053_ _12053_/A _12053_/B _12053_/C vssd1 vssd1 vccd1 vccd1 _12054_/A sky130_fd_sc_hd__and3_1
XFILLER_77_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11004_ _11004_/A vssd1 vssd1 vccd1 vccd1 _15614_/D sky130_fd_sc_hd__clkbuf_1
X_15812_ _07603_/A _15812_/D vssd1 vssd1 vccd1 vccd1 _15812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_15743_ _15763_/CLK _15743_/D vssd1 vssd1 vccd1 vccd1 _15743_/Q sky130_fd_sc_hd__dfxtp_1
X_12955_ _15923_/Q _12962_/C _07672_/A vssd1 vssd1 vccd1 vccd1 _12955_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11906_ _15763_/Q _15762_/Q _15761_/Q _11847_/X vssd1 vssd1 vccd1 vccd1 _15755_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15683_/CLK _15674_/D vssd1 vssd1 vccd1 vccd1 _15674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12886_ _12886_/A vssd1 vssd1 vccd1 vccd1 _15910_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _13250_/A vssd1 vssd1 vccd1 vccd1 _12972_/A sky130_fd_sc_hd__clkbuf_2
X_14625_ _16238_/Q _14778_/B _14627_/C vssd1 vssd1 vccd1 vccd1 _14630_/A sky130_fd_sc_hd__and3_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14561_/A _14555_/Y _14551_/B _14552_/C vssd1 vssd1 vccd1 vccd1 _14558_/B
+ sky130_fd_sc_hd__o211a_1
X_11768_ _15735_/Q _11774_/C _11713_/X vssd1 vssd1 vccd1 vccd1 _11768_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10719_ _10719_/A vssd1 vssd1 vccd1 vccd1 _15569_/D sky130_fd_sc_hd__clkbuf_1
X_13507_ _13507_/A _13507_/B vssd1 vssd1 vccd1 vccd1 _13509_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ _16205_/Q _14486_/C _07674_/A vssd1 vssd1 vccd1 vccd1 _14488_/B sky130_fd_sc_hd__a21o_1
X_11699_ _11697_/Y _11693_/C _11695_/X _11696_/Y vssd1 vssd1 vccd1 vccd1 _11700_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16226_ _16241_/CLK _16226_/D vssd1 vssd1 vccd1 vccd1 _16226_/Q sky130_fd_sc_hd__dfxtp_2
X_13438_ _16005_/Q _13445_/C _13437_/X vssd1 vssd1 vccd1 vccd1 _13438_/Y sky130_fd_sc_hd__a21oi_1
X_16157_ _16166_/CLK _16157_/D vssd1 vssd1 vccd1 vccd1 _16157_/Q sky130_fd_sc_hd__dfxtp_1
X_13369_ _13380_/C vssd1 vssd1 vccd1 vccd1 _13394_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ _16349_/Q _15107_/C _13950_/B vssd1 vssd1 vccd1 vccd1 _15109_/B sky130_fd_sc_hd__a21oi_1
X_16088_ _16367_/CLK _16088_/D vssd1 vssd1 vccd1 vccd1 _16088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07930_ _07930_/A _07930_/B vssd1 vssd1 vccd1 vccd1 _07932_/B sky130_fd_sc_hd__xor2_1
X_15039_ _15039_/A _15039_/B vssd1 vssd1 vccd1 vccd1 _15040_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07861_ _12077_/A _07861_/B vssd1 vssd1 vccd1 vccd1 _07887_/A sky130_fd_sc_hd__xnor2_4
XFILLER_122_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09600_ _15403_/Q _15402_/Q _15401_/Q _09541_/X vssd1 vssd1 vccd1 vccd1 _15395_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07792_ _16206_/Q vssd1 vssd1 vccd1 vccd1 _14546_/C sky130_fd_sc_hd__clkinv_4
XFILLER_37_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09531_ _09531_/A _09531_/B vssd1 vssd1 vccd1 vccd1 _09533_/B sky130_fd_sc_hd__nor2_1
X_09462_ _15374_/Q _09524_/B _09466_/C vssd1 vssd1 vccd1 vccd1 _09462_/Y sky130_fd_sc_hd__nand3_1
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08413_ _08413_/A vssd1 vssd1 vccd1 vccd1 _15212_/D sky130_fd_sc_hd__clkbuf_1
X_09393_ _09391_/Y _09384_/C _09386_/X _09387_/Y vssd1 vssd1 vccd1 vccd1 _09394_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08344_ _08344_/A _08344_/B vssd1 vssd1 vccd1 vccd1 _08384_/B sky130_fd_sc_hd__or2_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08275_ _15208_/Q _08279_/A _08429_/C vssd1 vssd1 vccd1 vccd1 _08275_/X sky130_fd_sc_hd__and3_1
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _09727_/X _09728_/Y _09724_/B _09725_/C vssd1 vssd1 vccd1 vccd1 _09731_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_43_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12740_ _12740_/A _12740_/B _12740_/C vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__and3_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12667_/X _12669_/Y _12670_/Y _12665_/C vssd1 vssd1 vccd1 vccd1 _12673_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14532_/A _14410_/B vssd1 vssd1 vccd1 vccd1 _14411_/B sky130_fd_sc_hd__and2_1
X_11622_ _11643_/C vssd1 vssd1 vccd1 vccd1 _11655_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15390_ _15484_/CLK _15390_/D vssd1 vssd1 vccd1 vccd1 _15390_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14341_ _14342_/B _14342_/C _14342_/A vssd1 vssd1 vccd1 vccd1 _14343_/B sky130_fd_sc_hd__a21o_1
XFILLER_11_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11553_ _11780_/A _11556_/C vssd1 vssd1 vccd1 vccd1 _11553_/X sky130_fd_sc_hd__or2_1
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10504_ _10504_/A vssd1 vssd1 vccd1 vccd1 _15535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14272_ _14269_/X _14272_/B vssd1 vssd1 vccd1 vccd1 _14272_/X sky130_fd_sc_hd__and2b_1
X_11484_ _11509_/A _11484_/B _11491_/B vssd1 vssd1 vccd1 vccd1 _15689_/D sky130_fd_sc_hd__nor3_1
X_16011_ _16011_/CLK _16011_/D vssd1 vssd1 vccd1 vccd1 _16011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13223_ _13223_/A _13223_/B _13223_/C vssd1 vssd1 vccd1 vccd1 _13224_/A sky130_fd_sc_hd__and3_1
X_10435_ _10432_/X _10433_/Y _10434_/Y _10430_/C vssd1 vssd1 vccd1 vccd1 _10437_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_137_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ _13617_/A vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__buf_2
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10366_ _10363_/X _10365_/Y _10360_/B _10361_/C vssd1 vssd1 vccd1 vccd1 _10368_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_88_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12112_/A _12105_/B _12105_/C vssd1 vssd1 vccd1 vccd1 _12106_/A sky130_fd_sc_hd__and3_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13283_/A vssd1 vssd1 vccd1 vccd1 _13149_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10297_ _10353_/A _10297_/B _10301_/A vssd1 vssd1 vccd1 vccd1 _15504_/D sky130_fd_sc_hd__nor3_1
XFILLER_88_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12036_ _12030_/B _12031_/C _12033_/X _12034_/Y vssd1 vssd1 vccd1 vccd1 _12037_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13987_ _13987_/A vssd1 vssd1 vccd1 vccd1 _16100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15726_ _15763_/CLK _15726_/D vssd1 vssd1 vccd1 vccd1 _15726_/Q sky130_fd_sc_hd__dfxtp_1
X_12938_ _12938_/A _12938_/B _12938_/C vssd1 vssd1 vccd1 vccd1 _12939_/C sky130_fd_sc_hd__nand3_1
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15657_ _15763_/CLK _15657_/D vssd1 vssd1 vccd1 vccd1 _15657_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12869_/A _12869_/B _12869_/C vssd1 vssd1 vccd1 vccd1 _12871_/B sky130_fd_sc_hd__or3_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ _14604_/Y _14607_/X _14528_/X vssd1 vssd1 vccd1 vccd1 _14608_/Y sky130_fd_sc_hd__a21oi_1
X_15588_ _15194_/Q _15588_/D vssd1 vssd1 vccd1 vccd1 _15588_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14539_ _14539_/A _14539_/B vssd1 vssd1 vccd1 vccd1 _16214_/D sky130_fd_sc_hd__nor2_1
XFILLER_147_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08060_ _07818_/A _07818_/B _08059_/X vssd1 vssd1 vccd1 vccd1 _08062_/B sky130_fd_sc_hd__o21a_1
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16209_ _16240_/CLK _16209_/D vssd1 vssd1 vccd1 vccd1 _16209_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ _08961_/B _08961_/C _08726_/X vssd1 vssd1 vccd1 vccd1 _08963_/C sky130_fd_sc_hd__o21ai_1
XFILLER_142_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07913_ _16323_/Q vssd1 vssd1 vccd1 vccd1 _07960_/A sky130_fd_sc_hd__inv_2
X_08893_ _08893_/A _08897_/C vssd1 vssd1 vccd1 vccd1 _08893_/X sky130_fd_sc_hd__or2_1
XFILLER_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07844_ _07844_/A _07844_/B vssd1 vssd1 vccd1 vccd1 _08022_/B sky130_fd_sc_hd__xor2_4
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07775_ _15575_/Q _08088_/B vssd1 vssd1 vccd1 vccd1 _07778_/B sky130_fd_sc_hd__xnor2_2
XFILLER_25_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09514_ _15383_/Q _09740_/B _09522_/C vssd1 vssd1 vccd1 vccd1 _09514_/X sky130_fd_sc_hd__and3_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09445_ _15373_/Q _09446_/C _09220_/X vssd1 vssd1 vccd1 vccd1 _09445_/Y sky130_fd_sc_hd__a21oi_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _09377_/B _09377_/C _09377_/A vssd1 vssd1 vccd1 vccd1 _09378_/B sky130_fd_sc_hd__a21o_1
X_08327_ _08365_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08329_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08258_ _08318_/A _08318_/B vssd1 vssd1 vccd1 vccd1 _08259_/B sky130_fd_sc_hd__xor2_4
XFILLER_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08189_ _07975_/A _07975_/B _07974_/A vssd1 vssd1 vccd1 vccd1 _08191_/C sky130_fd_sc_hd__a21oi_1
XFILLER_146_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10220_ _15493_/Q _10220_/B _10220_/C vssd1 vssd1 vccd1 vccd1 _10228_/B sky130_fd_sc_hd__and3_1
XFILLER_133_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _10148_/X _10149_/Y _10150_/Y _10146_/C vssd1 vssd1 vccd1 vccd1 _10153_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10082_ _15472_/Q _10310_/B _10085_/C vssd1 vssd1 vccd1 vccd1 _10082_/X sky130_fd_sc_hd__and3_1
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13910_ _15005_/A vssd1 vssd1 vccd1 vccd1 _15189_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14890_ _15005_/A vssd1 vssd1 vccd1 vccd1 _15051_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13841_ _16076_/Q _14088_/B _13846_/C vssd1 vssd1 vccd1 vccd1 _13841_/Y sky130_fd_sc_hd__nand3_1
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13772_ _16079_/Q _16078_/Q _16077_/Q _13723_/X vssd1 vssd1 vccd1 vccd1 _16062_/D
+ sky130_fd_sc_hd__o31a_1
X_10984_ _15619_/Q _15618_/Q _15617_/Q _10983_/X vssd1 vssd1 vccd1 vccd1 _15611_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15511_ _15224_/Q _15511_/D vssd1 vssd1 vccd1 vccd1 _15511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12723_ _12717_/B _12718_/C _12720_/X _12721_/Y vssd1 vssd1 vccd1 vccd1 _12724_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15442_ _15483_/CLK _15442_/D vssd1 vssd1 vccd1 vccd1 _15442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12654_ _12654_/A vssd1 vssd1 vccd1 vccd1 _12654_/X sky130_fd_sc_hd__buf_2
X_11605_ _15709_/Q _11719_/B _11605_/C vssd1 vssd1 vccd1 vccd1 _11614_/B sky130_fd_sc_hd__and3_1
X_15373_ _15484_/CLK _15373_/D vssd1 vssd1 vccd1 vccd1 _15373_/Q sky130_fd_sc_hd__dfxtp_1
X_12585_ _12621_/A _12585_/B _12585_/C vssd1 vssd1 vccd1 vccd1 _12586_/A sky130_fd_sc_hd__and3_1
X_11536_ _11533_/X _11534_/Y _11535_/Y _11531_/C vssd1 vssd1 vccd1 vccd1 _11538_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_11_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14324_ _14195_/X _14321_/B _14323_/Y vssd1 vssd1 vccd1 vccd1 _16168_/D sky130_fd_sc_hd__o21a_1
X_14255_ _14255_/A vssd1 vssd1 vccd1 vccd1 _16154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11467_ _11463_/X _11464_/Y _11466_/Y _11461_/C vssd1 vssd1 vccd1 vccd1 _11469_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _15086_/A vssd1 vssd1 vccd1 vccd1 _13206_/X sky130_fd_sc_hd__clkbuf_2
X_10418_ _15524_/Q _10590_/B _10426_/C vssd1 vssd1 vccd1 vccd1 _10421_/B sky130_fd_sc_hd__nand3_1
XFILLER_124_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14186_ _16142_/Q _14185_/C _14004_/X vssd1 vssd1 vccd1 vccd1 _14187_/B sky130_fd_sc_hd__a21o_1
X_11398_ _11398_/A _11398_/B _11398_/C vssd1 vssd1 vccd1 vccd1 _11399_/C sky130_fd_sc_hd__nand3_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _13654_/A vssd1 vssd1 vccd1 vccd1 _13349_/B sky130_fd_sc_hd__clkbuf_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _10375_/C vssd1 vssd1 vccd1 vccd1 _10389_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13066_/Y _13062_/C _13064_/X _13065_/Y vssd1 vssd1 vccd1 vccd1 _13069_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12019_ _15779_/Q _15781_/Q _15780_/Q _11847_/X vssd1 vssd1 vccd1 vccd1 _15773_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15709_ _15763_/CLK _15709_/D vssd1 vssd1 vccd1 vccd1 _15709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09230_ _15338_/Q _09285_/B _09236_/C vssd1 vssd1 vccd1 vccd1 _09230_/Y sky130_fd_sc_hd__nand3_1
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ _09158_/X _09159_/Y _09160_/Y _09156_/C vssd1 vssd1 vccd1 vccd1 _09163_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08112_ _15377_/Q vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__inv_2
X_09092_ _09093_/B _09093_/C _09093_/A vssd1 vssd1 vccd1 vccd1 _09094_/B sky130_fd_sc_hd__a21o_1
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08043_ _08043_/A _08182_/A vssd1 vssd1 vccd1 vccd1 _08147_/A sky130_fd_sc_hd__xnor2_4
XFILLER_107_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09994_ _10049_/A _09997_/C vssd1 vssd1 vccd1 vccd1 _09994_/X sky130_fd_sc_hd__or2_1
X_08945_ _15295_/Q _09001_/B _08945_/C vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__and3_1
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08876_ _08872_/X _08874_/Y _08875_/Y _08870_/C vssd1 vssd1 vccd1 vccd1 _08878_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_130_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07827_ _10347_/A _07827_/B vssd1 vssd1 vccd1 vccd1 _07828_/B sky130_fd_sc_hd__xnor2_4
XFILLER_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07758_ _15548_/Q _08140_/B vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__xnor2_4
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07689_ _08722_/A vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__buf_2
XFILLER_25_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09428_ _15370_/Q _09466_/C _09316_/X vssd1 vssd1 vccd1 vccd1 _09431_/B sky130_fd_sc_hd__a21oi_1
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09359_ _09472_/A _09362_/C vssd1 vssd1 vccd1 vccd1 _09359_/X sky130_fd_sc_hd__or2_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12370_ _12654_/A vssd1 vssd1 vccd1 vccd1 _12370_/X sky130_fd_sc_hd__buf_2
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11321_ _11321_/A _11321_/B vssd1 vssd1 vccd1 vccd1 _11326_/C sky130_fd_sc_hd__nor2_1
XFILLER_109_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14040_ _14040_/A _14040_/B vssd1 vssd1 vccd1 vccd1 _14040_/Y sky130_fd_sc_hd__nor2_1
X_11252_ _11826_/A vssd1 vssd1 vccd1 vccd1 _11373_/A sky130_fd_sc_hd__buf_2
XFILLER_109_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10203_ _10203_/A vssd1 vssd1 vccd1 vccd1 _15489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11183_ _15644_/Q _11244_/B _11191_/C vssd1 vssd1 vccd1 vccd1 _11183_/X sky130_fd_sc_hd__and3_1
XFILLER_69_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10134_ _10134_/A vssd1 vssd1 vccd1 vccd1 _10363_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15991_ _16007_/CLK _15991_/D vssd1 vssd1 vccd1 vccd1 _15991_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10065_ _10065_/A vssd1 vssd1 vccd1 vccd1 _10298_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14942_ _14980_/A vssd1 vssd1 vccd1 vccd1 _14942_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14873_ _14866_/B _14867_/C _14878_/A _14871_/Y vssd1 vssd1 vccd1 vccd1 _14878_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_29_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13824_ _16074_/Q _14071_/B _13824_/C vssd1 vssd1 vccd1 vccd1 _13829_/A sky130_fd_sc_hd__and3_1
XFILLER_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13755_ _13761_/A _13753_/Y _13754_/Y _13749_/C vssd1 vssd1 vccd1 vccd1 _13757_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10967_ _10965_/Y _10960_/C _10973_/A _10964_/Y vssd1 vssd1 vccd1 vccd1 _10973_/B
+ sky130_fd_sc_hd__a211oi_1
X_12706_ _12706_/A vssd1 vssd1 vccd1 vccd1 _12720_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13686_ _16049_/Q _13738_/B _13686_/C vssd1 vssd1 vccd1 vccd1 _13686_/X sky130_fd_sc_hd__and3_1
X_10898_ _15599_/Q _10904_/C _10897_/X vssd1 vssd1 vccd1 vccd1 _10898_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15425_ _15483_/CLK _15425_/D vssd1 vssd1 vccd1 vccd1 _15425_/Q sky130_fd_sc_hd__dfxtp_1
X_12637_ _12635_/A _12635_/B _12636_/X vssd1 vssd1 vccd1 vccd1 _15870_/D sky130_fd_sc_hd__a21oi_1
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15356_ _15356_/CLK _15356_/D vssd1 vssd1 vccd1 vccd1 _15356_/Q sky130_fd_sc_hd__dfxtp_1
X_12568_ _15861_/Q _12798_/B _12568_/C vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__and3_1
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14307_ _14307_/A _14307_/B vssd1 vssd1 vccd1 vccd1 _14307_/Y sky130_fd_sc_hd__nor2_1
X_11519_ _12377_/A vssd1 vssd1 vccd1 vccd1 _11519_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15287_ _15359_/CLK _15287_/D vssd1 vssd1 vccd1 vccd1 _15287_/Q sky130_fd_sc_hd__dfxtp_1
X_12499_ _15850_/Q _12500_/C _12384_/X vssd1 vssd1 vccd1 vccd1 _12499_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_144_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14238_ _14195_/X _14235_/B _14237_/Y vssd1 vssd1 vccd1 vccd1 _16150_/D sky130_fd_sc_hd__o21a_1
XFILLER_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14169_ _14343_/A _14169_/B _14169_/C vssd1 vssd1 vccd1 vccd1 _14170_/A sky130_fd_sc_hd__and3_1
XFILLER_124_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08730_ _15278_/Q _15277_/Q _15276_/Q _08604_/X vssd1 vssd1 vccd1 vccd1 _15261_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08661_ _13250_/A vssd1 vssd1 vccd1 vccd1 _14541_/A sky130_fd_sc_hd__buf_6
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07612_ _14414_/A vssd1 vssd1 vccd1 vccd1 _15030_/A sky130_fd_sc_hd__buf_4
XFILLER_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08592_ _08600_/B _08592_/B vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__or2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ _15337_/Q _09222_/C _09212_/X vssd1 vssd1 vccd1 vccd1 _09213_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09144_ _15326_/Q _09372_/B _09152_/C vssd1 vssd1 vccd1 vccd1 _09149_/A sky130_fd_sc_hd__and3_1
X_09075_ _09133_/A _09075_/B _09075_/C vssd1 vssd1 vccd1 vccd1 _09077_/B sky130_fd_sc_hd__or3_1
XFILLER_147_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08026_ _07844_/A _07844_/B _08025_/X vssd1 vssd1 vccd1 vccd1 _08035_/A sky130_fd_sc_hd__o21ai_4
XFILLER_107_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09977_ _09977_/A _09977_/B _09977_/C vssd1 vssd1 vccd1 vccd1 _09978_/A sky130_fd_sc_hd__and3_1
XFILLER_130_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08928_ _15293_/Q _09158_/B _08931_/C vssd1 vssd1 vccd1 vccd1 _08928_/X sky130_fd_sc_hd__and3_1
X_08859_ _15283_/Q _08919_/B _08859_/C vssd1 vssd1 vccd1 vccd1 _08859_/X sky130_fd_sc_hd__and3_1
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11870_ _15751_/Q _12099_/B _11872_/C vssd1 vssd1 vccd1 vccd1 _11870_/X sky130_fd_sc_hd__and3_1
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10821_ _10822_/B _10822_/C _10822_/A vssd1 vssd1 vccd1 vccd1 _10823_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10752_ _10750_/B _10750_/C _10751_/X vssd1 vssd1 vccd1 vccd1 _10753_/C sky130_fd_sc_hd__o21ai_1
XFILLER_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13540_ _13612_/A vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _13484_/C vssd1 vssd1 vccd1 vccd1 _13498_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10683_ _10681_/Y _10676_/C _10688_/A _10680_/Y vssd1 vssd1 vccd1 vccd1 _10688_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15210_ _16224_/CLK _15210_/D vssd1 vssd1 vccd1 vccd1 _15210_/Q sky130_fd_sc_hd__dfxtp_1
X_12422_ _12443_/C vssd1 vssd1 vccd1 vccd1 _12456_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16190_ _16247_/CLK _16190_/D vssd1 vssd1 vccd1 vccd1 _16190_/Q sky130_fd_sc_hd__dfxtp_2
X_15141_ _15175_/A _15141_/B _15145_/B vssd1 vssd1 vccd1 vccd1 _16353_/D sky130_fd_sc_hd__nor3_1
X_12353_ _12351_/A _12351_/B _12352_/X vssd1 vssd1 vccd1 vccd1 _15825_/D sky130_fd_sc_hd__a21oi_1
XFILLER_139_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11304_ _15662_/Q _11533_/B _11311_/C vssd1 vssd1 vccd1 vccd1 _11304_/X sky130_fd_sc_hd__and3_1
X_15072_ hold15/X _15142_/B _15072_/C vssd1 vssd1 vccd1 vccd1 _15074_/A sky130_fd_sc_hd__and3_1
X_12284_ _15816_/Q _12512_/B _12284_/C vssd1 vssd1 vccd1 vccd1 _12294_/A sky130_fd_sc_hd__and3_1
XFILLER_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14023_ _14098_/A _14023_/B _14028_/A vssd1 vssd1 vccd1 vccd1 _16108_/D sky130_fd_sc_hd__nor3_1
X_11235_ _11235_/A vssd1 vssd1 vccd1 vccd1 _15650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11166_ _11166_/A _11166_/B _11166_/C vssd1 vssd1 vccd1 vccd1 _11167_/C sky130_fd_sc_hd__nand3_1
XFILLER_95_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10117_ _10153_/A _10117_/B _10117_/C vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__and3_1
XFILLER_110_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11097_ _11097_/A vssd1 vssd1 vccd1 vccd1 _15628_/D sky130_fd_sc_hd__clkbuf_1
X_15974_ _15984_/CLK _15974_/D vssd1 vssd1 vccd1 vccd1 _15974_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10048_ _10048_/A _10048_/B vssd1 vssd1 vccd1 vccd1 _10053_/C sky130_fd_sc_hd__nor2_1
X_14925_ _15045_/A _14930_/C vssd1 vssd1 vccd1 vccd1 _14925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14856_ _14772_/X _14855_/A _14815_/X vssd1 vssd1 vccd1 vccd1 _14856_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13807_ _13812_/B _13807_/B vssd1 vssd1 vccd1 vccd1 _13809_/A sky130_fd_sc_hd__or2_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14787_ _14787_/A vssd1 vssd1 vccd1 vccd1 _16271_/D sky130_fd_sc_hd__clkbuf_1
X_11999_ _12853_/A vssd1 vssd1 vccd1 vccd1 _12228_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13738_ _16058_/Q _13738_/B _13738_/C vssd1 vssd1 vccd1 vccd1 _13738_/X sky130_fd_sc_hd__and3_1
X_13669_ _16061_/Q _16060_/Q _16059_/Q _13467_/X vssd1 vssd1 vccd1 vccd1 _16044_/D
+ sky130_fd_sc_hd__o31a_1
X_15408_ _15483_/CLK _15408_/D vssd1 vssd1 vccd1 vccd1 _15408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15339_ _15339_/CLK _15339_/D vssd1 vssd1 vccd1 vccd1 _15339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09900_ _09900_/A _09900_/B _09900_/C vssd1 vssd1 vccd1 vccd1 _09901_/C sky130_fd_sc_hd__nand3_1
XFILLER_59_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _10983_/A vssd1 vssd1 vccd1 vccd1 _09831_/X sky130_fd_sc_hd__clkbuf_2
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09762_ _09825_/A vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08711_/Y _08704_/C _08718_/A _08707_/Y vssd1 vssd1 vccd1 vccd1 _08718_/B
+ sky130_fd_sc_hd__a211oi_1
X_09693_ _09693_/A vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__buf_2
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08644_ _15249_/Q _08651_/C _08575_/X vssd1 vssd1 vccd1 vccd1 _08644_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08575_ _13064_/B vssd1 vssd1 vccd1 vccd1 _08575_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09127_ _09133_/B _09127_/B vssd1 vssd1 vccd1 vccd1 _09129_/A sky130_fd_sc_hd__or2_1
XFILLER_135_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09058_ _09058_/A _09058_/B _09058_/C vssd1 vssd1 vccd1 vccd1 _09059_/A sky130_fd_sc_hd__and3_1
XFILLER_135_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08009_ _08010_/A _08010_/B vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11020_ _11020_/A vssd1 vssd1 vccd1 vccd1 _15616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12971_ _12971_/A _12971_/B vssd1 vssd1 vccd1 vccd1 _12973_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14710_ _14748_/A _14710_/B _14710_/C vssd1 vssd1 vccd1 vccd1 _14711_/A sky130_fd_sc_hd__and3_1
X_11922_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15690_ _15763_/CLK _15690_/D vssd1 vssd1 vccd1 vccd1 _15690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14641_ _14641_/A _14641_/B vssd1 vssd1 vccd1 vccd1 _14643_/A sky130_fd_sc_hd__or2_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11853_ _15748_/Q _11891_/C _11624_/X vssd1 vssd1 vccd1 vccd1 _11855_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10804_ _10802_/A _10802_/B _10803_/X vssd1 vssd1 vccd1 vccd1 _15582_/D sky130_fd_sc_hd__a21oi_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11784_ _12015_/A _11784_/B _11784_/C vssd1 vssd1 vccd1 vccd1 _11786_/B sky130_fd_sc_hd__or3_1
X_14572_ _14806_/A _14572_/B vssd1 vssd1 vccd1 vccd1 _14573_/B sky130_fd_sc_hd__and2_1
X_16311_ _16317_/CLK _16311_/D vssd1 vssd1 vccd1 vccd1 _16311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13523_ _16020_/Q _13675_/B _13523_/C vssd1 vssd1 vccd1 vccd1 _13529_/A sky130_fd_sc_hd__and3_1
X_10735_ _15573_/Q _10741_/C _10562_/X vssd1 vssd1 vccd1 vccd1 _10735_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16242_ _16242_/CLK hold25/X vssd1 vssd1 vccd1 vccd1 _16242_/Q sky130_fd_sc_hd__dfxtp_1
X_10666_ _10662_/X _10664_/Y _10665_/Y _10659_/C vssd1 vssd1 vccd1 vccd1 _10668_/B
+ sky130_fd_sc_hd__o211ai_1
X_13454_ _13460_/B _13454_/B vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__or2_1
XFILLER_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12405_ _15835_/Q _12575_/B _12405_/C vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__and3_1
X_16173_ _16192_/CLK _16173_/D vssd1 vssd1 vccd1 vccd1 _16173_/Q sky130_fd_sc_hd__dfxtp_2
X_13385_ _13385_/A vssd1 vssd1 vccd1 vccd1 _15993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10597_ _15552_/Q _10604_/C _10364_/X vssd1 vssd1 vccd1 vccd1 _10597_/Y sky130_fd_sc_hd__a21oi_1
X_15124_ _15013_/X _15122_/A _15123_/Y vssd1 vssd1 vccd1 vccd1 _16349_/D sky130_fd_sc_hd__o21a_1
X_12336_ _12334_/Y _12329_/C _12331_/X _12333_/Y vssd1 vssd1 vccd1 vccd1 _12337_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12267_ _12267_/A vssd1 vssd1 vccd1 vccd1 _15812_/D sky130_fd_sc_hd__clkbuf_1
X_15055_ _15013_/X _15053_/A _15054_/Y vssd1 vssd1 vccd1 vccd1 _16331_/D sky130_fd_sc_hd__o21a_1
XFILLER_126_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11218_ _11507_/A vssd1 vssd1 vccd1 vccd1 _11449_/B sky130_fd_sc_hd__buf_2
X_14006_ _14003_/X _14006_/B vssd1 vssd1 vccd1 vccd1 _14006_/X sky130_fd_sc_hd__and2b_1
X_12198_ _15802_/Q _12235_/C _12197_/X vssd1 vssd1 vccd1 vccd1 _12200_/B sky130_fd_sc_hd__a21oi_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11149_ _11147_/A _11147_/B _11148_/X vssd1 vssd1 vccd1 vccd1 _15636_/D sky130_fd_sc_hd__a21oi_1
XFILLER_83_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15957_ _15970_/CLK _15957_/D vssd1 vssd1 vccd1 vccd1 _15957_/Q sky130_fd_sc_hd__dfxtp_1
X_14908_ _14908_/A _14908_/B _14908_/C vssd1 vssd1 vccd1 vccd1 _14909_/C sky130_fd_sc_hd__nand3_1
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15888_ _07603_/A _15888_/D vssd1 vssd1 vccd1 vccd1 _15888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14839_ _16286_/Q _14838_/C _14718_/X vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08360_ _08321_/A _08321_/B _08359_/Y vssd1 vssd1 vccd1 vccd1 _08381_/B sky130_fd_sc_hd__a21oi_2
XFILLER_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08291_ _08291_/A _08193_/A vssd1 vssd1 vccd1 vccd1 _08293_/A sky130_fd_sc_hd__or2b_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09814_ _09820_/A _09812_/Y _09813_/Y _09807_/C vssd1 vssd1 vccd1 vccd1 _09816_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09745_ _09743_/Y _09738_/C _09740_/X _09742_/Y vssd1 vssd1 vccd1 vccd1 _09746_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09676_/A vssd1 vssd1 vccd1 vccd1 _15407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _08622_/X _08626_/Y _08619_/B _08620_/C vssd1 vssd1 vccd1 vccd1 _08629_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08558_ _08580_/A hold35/X _08558_/C vssd1 vssd1 vccd1 vccd1 _08559_/A sky130_fd_sc_hd__and3_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08489_ _08519_/A _08489_/B _08489_/C vssd1 vssd1 vccd1 vccd1 _08490_/A sky130_fd_sc_hd__and3_1
XFILLER_23_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10520_ _10577_/A _10520_/B _10520_/C vssd1 vssd1 vccd1 vccd1 _10522_/B sky130_fd_sc_hd__or3_1
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _10449_/Y _10444_/C _10456_/A _10447_/Y vssd1 vssd1 vccd1 vccd1 _10456_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_109_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13170_ _13223_/A _13170_/B _13170_/C vssd1 vssd1 vccd1 vccd1 _13171_/A sky130_fd_sc_hd__and3_1
XFILLER_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10382_ _15518_/Q _10389_/C _10318_/X vssd1 vssd1 vccd1 vccd1 _10382_/Y sky130_fd_sc_hd__a21oi_1
X_12121_ _15790_/Q _12291_/B _12121_/C vssd1 vssd1 vccd1 vccd1 _12130_/B sky130_fd_sc_hd__and3_1
XFILLER_124_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12052_ _12050_/Y _12045_/C _12047_/X _12049_/Y vssd1 vssd1 vccd1 vccd1 _12053_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11003_ _11019_/A _11003_/B _11003_/C vssd1 vssd1 vccd1 vccd1 _11004_/A sky130_fd_sc_hd__and3_1
XFILLER_77_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15811_ _07603_/A _15811_/D vssd1 vssd1 vccd1 vccd1 _15811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15742_ _15794_/CLK _15742_/D vssd1 vssd1 vccd1 vccd1 _15742_/Q sky130_fd_sc_hd__dfxtp_1
X_12954_ _15923_/Q _12954_/B _12962_/C vssd1 vssd1 vccd1 vccd1 _12954_/X sky130_fd_sc_hd__and3_1
XFILLER_18_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11905_ _11905_/A vssd1 vssd1 vccd1 vccd1 _15754_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _15763_/CLK _15673_/D vssd1 vssd1 vccd1 vccd1 _15673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _12906_/A _12885_/B _12885_/C vssd1 vssd1 vccd1 vccd1 _12886_/A sky130_fd_sc_hd__and3_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _15021_/A vssd1 vssd1 vccd1 vccd1 _14778_/B sky130_fd_sc_hd__buf_2
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11836_/A _11836_/B vssd1 vssd1 vccd1 vccd1 _11839_/B sky130_fd_sc_hd__nor2_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _16221_/Q _14554_/C _14634_/B vssd1 vssd1 vccd1 vccd1 _14555_/Y sky130_fd_sc_hd__a21oi_1
X_11767_ _15735_/Q _11943_/B _11767_/C vssd1 vssd1 vccd1 vccd1 _11778_/A sky130_fd_sc_hd__and3_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _13512_/B _13506_/B vssd1 vssd1 vccd1 vccd1 _13509_/A sky130_fd_sc_hd__or2_1
X_10718_ _10732_/A _10718_/B _10718_/C vssd1 vssd1 vccd1 vccd1 _10719_/A sky130_fd_sc_hd__and3_1
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ _16205_/Q _14566_/B _14486_/C vssd1 vssd1 vccd1 vccd1 _14486_/X sky130_fd_sc_hd__and3_1
XFILLER_146_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11698_ _11695_/X _11696_/Y _11697_/Y _11693_/C vssd1 vssd1 vccd1 vccd1 _11700_/B
+ sky130_fd_sc_hd__o211ai_1
X_16225_ _16359_/CLK _16225_/D vssd1 vssd1 vccd1 vccd1 _16225_/Q sky130_fd_sc_hd__dfxtp_2
X_13437_ _13693_/A vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_127_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10649_ _15560_/Q _10654_/C _10648_/X vssd1 vssd1 vccd1 vccd1 _10651_/C sky130_fd_sc_hd__a21o_1
X_16156_ _16166_/CLK _16156_/D vssd1 vssd1 vccd1 vccd1 _16156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13368_ _13372_/C vssd1 vssd1 vccd1 vccd1 _13380_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15107_ _16349_/Q _15142_/B _15107_/C vssd1 vssd1 vccd1 vccd1 _15109_/A sky130_fd_sc_hd__and3_1
X_12319_ _12317_/X _12318_/Y _12314_/B _12315_/C vssd1 vssd1 vccd1 vccd1 _12321_/B
+ sky130_fd_sc_hd__o211ai_1
X_16087_ _16367_/CLK _16087_/D vssd1 vssd1 vccd1 vccd1 _16087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13299_ _13304_/B _13299_/B vssd1 vssd1 vccd1 vccd1 _13301_/A sky130_fd_sc_hd__or2_1
X_15038_ _15038_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _15040_/A sky130_fd_sc_hd__or2_1
XFILLER_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07860_ _07860_/A _07860_/B vssd1 vssd1 vccd1 vccd1 _07861_/B sky130_fd_sc_hd__nand2_2
XFILLER_95_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07791_ _15908_/Q vssd1 vssd1 vccd1 vccd1 _12874_/A sky130_fd_sc_hd__inv_2
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ _09537_/B _09530_/B vssd1 vssd1 vccd1 vccd1 _09533_/A sky130_fd_sc_hd__or2_1
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09461_ _15375_/Q _09466_/C _09404_/X vssd1 vssd1 vccd1 vccd1 _09461_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08412_ _15017_/A _08412_/B _08412_/C vssd1 vssd1 vccd1 vccd1 _08413_/A sky130_fd_sc_hd__and3_1
X_09392_ _09386_/X _09387_/Y _09391_/Y _09384_/C vssd1 vssd1 vccd1 vccd1 _09394_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_52_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08343_ _08343_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ _08436_/A _08332_/B vssd1 vssd1 vccd1 vccd1 _08274_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07989_ _13824_/C _07989_/B vssd1 vssd1 vccd1 vccd1 _07989_/X sky130_fd_sc_hd__or2_1
X_09728_ _15417_/Q _09735_/C _09497_/X vssd1 vssd1 vccd1 vccd1 _09728_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09659_ _09671_/C vssd1 vssd1 vccd1 vccd1 _09680_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _15876_/Q _12840_/B _12670_/C vssd1 vssd1 vccd1 vccd1 _12670_/Y sky130_fd_sc_hd__nand3_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11635_/C vssd1 vssd1 vccd1 vccd1 _11643_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14340_ _16175_/Q _14345_/C _14250_/X vssd1 vssd1 vccd1 vccd1 _14342_/C sky130_fd_sc_hd__a21o_1
X_11552_ _11552_/A _11552_/B vssd1 vssd1 vccd1 vccd1 _11556_/C sky130_fd_sc_hd__nor2_1
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ _10503_/A _10503_/B _10503_/C vssd1 vssd1 vccd1 vccd1 _10504_/A sky130_fd_sc_hd__and3_1
XFILLER_128_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11483_ _11481_/Y _11477_/C _11491_/A _11480_/Y vssd1 vssd1 vccd1 vccd1 _11491_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_109_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14271_ _16160_/Q _14269_/C _14270_/X vssd1 vssd1 vccd1 vccd1 _14272_/B sky130_fd_sc_hd__a21o_1
X_16010_ _16011_/CLK _16010_/D vssd1 vssd1 vccd1 vccd1 _16010_/Q sky130_fd_sc_hd__dfxtp_2
X_10434_ _15525_/Q _10492_/B _10434_/C vssd1 vssd1 vccd1 vccd1 _10434_/Y sky130_fd_sc_hd__nand3_1
X_13222_ _13222_/A _13222_/B _13222_/C vssd1 vssd1 vccd1 vccd1 _13223_/C sky130_fd_sc_hd__nand3_1
X_10365_ _15516_/Q _10375_/C _10364_/X vssd1 vssd1 vccd1 vccd1 _10365_/Y sky130_fd_sc_hd__a21oi_1
X_13153_ _13666_/A vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__buf_2
XFILLER_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _12102_/Y _12097_/C _12099_/X _12101_/Y vssd1 vssd1 vccd1 vccd1 _12105_/C
+ sky130_fd_sc_hd__a211o_1
X_13084_ _13082_/A _13082_/B _13083_/X vssd1 vssd1 vccd1 vccd1 _15943_/D sky130_fd_sc_hd__a21oi_1
XFILLER_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10296_ _15505_/Q _10532_/B _10304_/C vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__and3_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12035_ _12033_/X _12034_/Y _12030_/B _12031_/C vssd1 vssd1 vccd1 vccd1 _12037_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_111_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13986_ _14029_/A _13986_/B _13986_/C vssd1 vssd1 vccd1 vccd1 _13987_/A sky130_fd_sc_hd__and3_1
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15725_ _15763_/CLK _15725_/D vssd1 vssd1 vccd1 vccd1 _15725_/Q sky130_fd_sc_hd__dfxtp_1
X_12937_ _12938_/B _12938_/C _12938_/A vssd1 vssd1 vccd1 vccd1 _12939_/B sky130_fd_sc_hd__a21o_1
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15656_ _15656_/CLK _15656_/D vssd1 vssd1 vccd1 vccd1 _15656_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12906_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14607_ _14605_/X _14607_/B vssd1 vssd1 vccd1 vccd1 _14607_/X sky130_fd_sc_hd__and2b_1
X_11819_ _15743_/Q _11819_/B _11827_/C vssd1 vssd1 vccd1 vccd1 _11819_/X sky130_fd_sc_hd__and3_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15587_ _15194_/Q _15587_/D vssd1 vssd1 vccd1 vccd1 _15587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _15897_/Q _12805_/C _12569_/X vssd1 vssd1 vccd1 vccd1 _12799_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14538_ _14368_/A _14372_/X _14533_/B _14459_/X vssd1 vssd1 vccd1 vccd1 _14539_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14469_ _16202_/Q _14474_/C _07632_/A vssd1 vssd1 vccd1 vccd1 _14471_/C sky130_fd_sc_hd__a21o_1
XFILLER_128_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16208_ _16247_/CLK _16208_/D vssd1 vssd1 vccd1 vccd1 _16208_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16139_ _16143_/CLK _16139_/D vssd1 vssd1 vccd1 vccd1 _16139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08961_ _09133_/A _08961_/B _08961_/C vssd1 vssd1 vccd1 vccd1 _08963_/B sky130_fd_sc_hd__or3_1
XFILLER_130_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07912_ _16008_/Q vssd1 vssd1 vccd1 vccd1 _13523_/C sky130_fd_sc_hd__clkinv_4
X_08892_ _08892_/A _08892_/B vssd1 vssd1 vccd1 vccd1 _08897_/C sky130_fd_sc_hd__nor2_1
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07843_ _13162_/C _07843_/B vssd1 vssd1 vccd1 vccd1 _07844_/B sky130_fd_sc_hd__xnor2_4
XFILLER_96_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07774_ _15557_/Q _15539_/Q vssd1 vssd1 vccd1 vccd1 _08088_/B sky130_fd_sc_hd__xor2_2
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09513_ _09801_/A vssd1 vssd1 vccd1 vccd1 _09740_/B sky130_fd_sc_hd__buf_2
XFILLER_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _15373_/Q _09444_/B _09446_/C vssd1 vssd1 vccd1 vccd1 _09444_/X sky130_fd_sc_hd__and3_1
XFILLER_25_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _15362_/Q _09380_/C _09205_/X vssd1 vssd1 vccd1 vccd1 _09377_/C sky130_fd_sc_hd__a21o_1
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08326_ _08338_/B _08326_/B vssd1 vssd1 vccd1 vccd1 _08328_/B sky130_fd_sc_hd__xor2_4
XFILLER_138_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08257_ _08143_/A _08143_/B _08256_/Y vssd1 vssd1 vccd1 vccd1 _08318_/B sky130_fd_sc_hd__a21oi_2
XFILLER_138_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_08188_ _08188_/A _08002_/A vssd1 vssd1 vccd1 vccd1 _08191_/B sky130_fd_sc_hd__or2b_1
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10150_ _15481_/Q _10150_/B _10155_/C vssd1 vssd1 vccd1 vccd1 _10150_/Y sky130_fd_sc_hd__nand3_1
X_10081_ _10081_/A vssd1 vssd1 vccd1 vccd1 _10310_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13840_ _14300_/A vssd1 vssd1 vccd1 vccd1 _14088_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13771_ _13666_/X _13768_/C _13770_/Y vssd1 vssd1 vccd1 vccd1 _16061_/D sky130_fd_sc_hd__a21oi_1
X_10983_ _10983_/A vssd1 vssd1 vccd1 vccd1 _10983_/X sky130_fd_sc_hd__buf_2
XFILLER_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15510_ _15224_/Q _15510_/D vssd1 vssd1 vccd1 vccd1 _15510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12722_ _12720_/X _12721_/Y _12717_/B _12718_/C vssd1 vssd1 vccd1 vccd1 _12724_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15441_ _15483_/CLK _15441_/D vssd1 vssd1 vccd1 vccd1 _15441_/Q sky130_fd_sc_hd__dfxtp_2
X_12653_ _15875_/Q _12653_/B _12660_/C vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__nand3_1
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11604_ _11661_/A _11604_/B _11608_/B vssd1 vssd1 vccd1 vccd1 _15707_/D sky130_fd_sc_hd__nor3_1
X_15372_ _15484_/CLK _15372_/D vssd1 vssd1 vccd1 vccd1 _15372_/Q sky130_fd_sc_hd__dfxtp_1
X_12584_ _12583_/B _12583_/C _12472_/X vssd1 vssd1 vccd1 vccd1 _12585_/C sky130_fd_sc_hd__o21ai_1
X_14323_ _14149_/X _14321_/B _14316_/X vssd1 vssd1 vccd1 vccd1 _14323_/Y sky130_fd_sc_hd__a21oi_1
X_11535_ _15697_/Q _11650_/B _11541_/C vssd1 vssd1 vccd1 vccd1 _11535_/Y sky130_fd_sc_hd__nand3_1
XFILLER_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14254_ _14343_/A _14254_/B _14254_/C vssd1 vssd1 vccd1 vccd1 _14255_/A sky130_fd_sc_hd__and3_1
X_11466_ _15687_/Q _11697_/B _11466_/C vssd1 vssd1 vccd1 vccd1 _11466_/Y sky130_fd_sc_hd__nand3_1
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ _13205_/A vssd1 vssd1 vccd1 vccd1 _15961_/D sky130_fd_sc_hd__clkbuf_1
X_10417_ _10511_/A _10417_/B _10421_/A vssd1 vssd1 vccd1 vccd1 _15522_/D sky130_fd_sc_hd__nor3_1
XFILLER_124_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11397_ _11398_/B _11398_/C _11398_/A vssd1 vssd1 vccd1 vccd1 _11399_/B sky130_fd_sc_hd__a21o_1
X_14185_ _16142_/Q _14357_/B _14185_/C vssd1 vssd1 vccd1 vccd1 _14185_/X sky130_fd_sc_hd__and3_1
X_13136_ _13218_/A _13136_/B _13141_/B vssd1 vssd1 vccd1 vccd1 _15950_/D sky130_fd_sc_hd__nor3_1
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _10363_/C vssd1 vssd1 vccd1 vccd1 _10375_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _10279_/A _10279_/B vssd1 vssd1 vccd1 vccd1 _10280_/B sky130_fd_sc_hd__nor2_1
X_13067_ _13064_/X _13065_/Y _13066_/Y _13062_/C vssd1 vssd1 vccd1 vccd1 _13069_/B
+ sky130_fd_sc_hd__o211ai_1
X_12018_ _12018_/A vssd1 vssd1 vccd1 vccd1 _15772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13969_ _14459_/A vssd1 vssd1 vccd1 vccd1 _13969_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15708_ _15763_/CLK _15708_/D vssd1 vssd1 vccd1 vccd1 _15708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15639_ _15655_/CLK _15639_/D vssd1 vssd1 vccd1 vccd1 _15639_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ _15328_/Q _09334_/B _09160_/C vssd1 vssd1 vccd1 vccd1 _09160_/Y sky130_fd_sc_hd__nand3_1
X_08111_ _15395_/Q vssd1 vssd1 vccd1 vccd1 _09601_/A sky130_fd_sc_hd__clkinv_2
XFILLER_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09091_ _15318_/Q _09096_/C _08913_/X vssd1 vssd1 vccd1 vccd1 _09093_/C sky130_fd_sc_hd__a21o_1
XFILLER_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08042_ _08042_/A _08042_/B vssd1 vssd1 vccd1 vccd1 _08182_/A sky130_fd_sc_hd__xnor2_2
XFILLER_134_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _09993_/A _09993_/B vssd1 vssd1 vccd1 vccd1 _09997_/C sky130_fd_sc_hd__nor2_1
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08944_ _08944_/A vssd1 vssd1 vccd1 vccd1 _09066_/A sky130_fd_sc_hd__buf_2
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08875_ _15284_/Q _08996_/B _08880_/C vssd1 vssd1 vccd1 vccd1 _08875_/Y sky130_fd_sc_hd__nand3_1
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07826_ _07826_/A _07826_/B vssd1 vssd1 vccd1 vccd1 _07827_/B sky130_fd_sc_hd__nand2_2
XFILLER_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07757_ _07757_/A _07757_/B vssd1 vssd1 vccd1 vccd1 _08140_/B sky130_fd_sc_hd__xor2_4
XFILLER_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07688_ _14964_/A vssd1 vssd1 vccd1 vccd1 _07688_/X sky130_fd_sc_hd__buf_2
XFILLER_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09427_ _09460_/C vssd1 vssd1 vccd1 vccd1 _09466_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09358_ _09358_/A _09358_/B vssd1 vssd1 vccd1 vccd1 _09362_/C sky130_fd_sc_hd__nor2_1
XFILLER_60_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08309_ _08251_/A _08251_/B _08250_/A vssd1 vssd1 vccd1 vccd1 _08384_/C sky130_fd_sc_hd__a21oi_1
XFILLER_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09289_ _09289_/A vssd1 vssd1 vccd1 vccd1 _15347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ _11320_/A _11320_/B vssd1 vssd1 vccd1 vccd1 _11321_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11251_ _11963_/A vssd1 vssd1 vccd1 vccd1 _11826_/A sky130_fd_sc_hd__buf_2
XFILLER_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ _10210_/A _10202_/B _10202_/C vssd1 vssd1 vccd1 vccd1 _10203_/A sky130_fd_sc_hd__and3_1
X_11182_ _11182_/A vssd1 vssd1 vccd1 vccd1 _15642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10133_ _10133_/A vssd1 vssd1 vccd1 vccd1 _15478_/D sky130_fd_sc_hd__clkbuf_1
X_15990_ _16007_/CLK _15990_/D vssd1 vssd1 vccd1 vccd1 _15990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10064_ _10064_/A _10064_/B _10071_/A vssd1 vssd1 vccd1 vccd1 _15468_/D sky130_fd_sc_hd__nor3_1
X_14941_ _16311_/Q _14941_/B _14941_/C vssd1 vssd1 vccd1 vccd1 _14945_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14872_ _14878_/A _14871_/Y _14866_/B _14867_/C vssd1 vssd1 vccd1 vccd1 _14874_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13823_ _16074_/Q _13853_/C _13822_/X vssd1 vssd1 vccd1 vccd1 _13825_/B sky130_fd_sc_hd__a21oi_1
XFILLER_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13754_ _16059_/Q _13801_/B _13758_/C vssd1 vssd1 vccd1 vccd1 _13754_/Y sky130_fd_sc_hd__nand3_1
X_10966_ _10973_/A _10964_/Y _10965_/Y _10960_/C vssd1 vssd1 vccd1 vccd1 _10968_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _15889_/Q _15888_/Q _15887_/Q _12704_/X vssd1 vssd1 vccd1 vccd1 _15881_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13685_ _13685_/A vssd1 vssd1 vccd1 vccd1 _16046_/D sky130_fd_sc_hd__clkbuf_1
X_10897_ _12048_/A vssd1 vssd1 vccd1 vccd1 _10897_/X sky130_fd_sc_hd__buf_2
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15424_ _15483_/CLK _15424_/D vssd1 vssd1 vccd1 vccd1 _15424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12636_ _12636_/A _12640_/C vssd1 vssd1 vccd1 vccd1 _12636_/X sky130_fd_sc_hd__or2_1
X_15355_ _15356_/CLK _15355_/D vssd1 vssd1 vccd1 vccd1 _15355_/Q sky130_fd_sc_hd__dfxtp_1
X_12567_ _12853_/A vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__clkbuf_2
X_14306_ _16168_/Q _14313_/C _14177_/X vssd1 vssd1 vccd1 vccd1 _14308_/B sky130_fd_sc_hd__a21oi_1
X_11518_ _15696_/Q _11576_/B _11518_/C vssd1 vssd1 vccd1 vccd1 _11518_/X sky130_fd_sc_hd__and3_1
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15286_ _15286_/CLK _15286_/D vssd1 vssd1 vccd1 vccd1 _15286_/Q sky130_fd_sc_hd__dfxtp_1
X_12498_ _15850_/Q _12667_/B _12500_/C vssd1 vssd1 vccd1 vccd1 _12498_/X sky130_fd_sc_hd__and3_1
XFILLER_144_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14237_ _14149_/X _14235_/B _14196_/X vssd1 vssd1 vccd1 vccd1 _14237_/Y sky130_fd_sc_hd__a21oi_1
X_11449_ _15685_/Q _11449_/B _11457_/C vssd1 vssd1 vccd1 vccd1 _11454_/A sky130_fd_sc_hd__and3_1
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14168_ _14168_/A _14168_/B _14168_/C vssd1 vssd1 vccd1 vccd1 _14169_/C sky130_fd_sc_hd__nand3_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13119_ _13532_/A vssd1 vssd1 vccd1 vccd1 _14080_/B sky130_fd_sc_hd__buf_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _16124_/Q _14099_/B _14099_/C vssd1 vssd1 vccd1 vccd1 _14106_/B sky130_fd_sc_hd__and3_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08660_ _08660_/A _08660_/B vssd1 vssd1 vccd1 vccd1 _08663_/B sky130_fd_sc_hd__nor2_1
XFILLER_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07611_ _13250_/A vssd1 vssd1 vccd1 vccd1 _14414_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08591_ _15242_/Q _08588_/C _08590_/X vssd1 vssd1 vccd1 vccd1 _08592_/B sky130_fd_sc_hd__a21oi_1
XFILLER_93_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ _13051_/B vssd1 vssd1 vccd1 vccd1 _09212_/X sky130_fd_sc_hd__buf_2
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09143_ _10007_/A vssd1 vssd1 vccd1 vccd1 _09372_/B sky130_fd_sc_hd__clkbuf_4
X_09074_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09115_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08025_ _14207_/C _08025_/B vssd1 vssd1 vccd1 vccd1 _08025_/X sky130_fd_sc_hd__or2_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09976_ _09974_/Y _09970_/C _09972_/X _09973_/Y vssd1 vssd1 vccd1 vccd1 _09977_/C
+ sky130_fd_sc_hd__a211o_1
X_08927_ _10081_/A vssd1 vssd1 vccd1 vccd1 _09158_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08858_ _08858_/A vssd1 vssd1 vccd1 vccd1 _15281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07809_ _16188_/Q vssd1 vssd1 vccd1 vccd1 _14466_/C sky130_fd_sc_hd__inv_6
X_08789_ _15261_/Q vssd1 vssd1 vccd1 vccd1 _08802_/C sky130_fd_sc_hd__clkinv_2
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10820_ _15587_/Q _10825_/C _10648_/X vssd1 vssd1 vccd1 vccd1 _10822_/C sky130_fd_sc_hd__a21o_1
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10751_ _10751_/A vssd1 vssd1 vccd1 vccd1 _10751_/X sky130_fd_sc_hd__buf_2
XFILLER_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13470_ _13475_/C vssd1 vssd1 vccd1 vccd1 _13484_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10682_ _10688_/A _10680_/Y _10681_/Y _10676_/C vssd1 vssd1 vccd1 vccd1 _10684_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12421_ _12434_/C vssd1 vssd1 vccd1 vccd1 _12443_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_138_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15140_ _15134_/B _15135_/C _15145_/A _15138_/Y vssd1 vssd1 vccd1 vccd1 _15145_/B
+ sky130_fd_sc_hd__a211oi_1
X_12352_ _12352_/A _12356_/C vssd1 vssd1 vccd1 vccd1 _12352_/X sky130_fd_sc_hd__or2_1
XFILLER_5_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11303_ _11303_/A vssd1 vssd1 vccd1 vccd1 _11533_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15071_ _15106_/A _15071_/B _15075_/B vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__nor3_1
X_12283_ _12853_/A vssd1 vssd1 vccd1 vccd1 _12512_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14022_ _16111_/Q _14117_/B _14022_/C vssd1 vssd1 vccd1 vccd1 _14028_/A sky130_fd_sc_hd__and3_1
X_11234_ _11249_/A _11234_/B _11234_/C vssd1 vssd1 vccd1 vccd1 _11235_/A sky130_fd_sc_hd__and3_1
XFILLER_106_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ _11166_/B _11166_/C _11166_/A vssd1 vssd1 vccd1 vccd1 _11167_/B sky130_fd_sc_hd__a21o_1
XFILLER_136_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10116_ _10115_/B _10115_/C _09884_/X vssd1 vssd1 vccd1 vccd1 _10117_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11096_ _11133_/A _11096_/B _11096_/C vssd1 vssd1 vccd1 vccd1 _11097_/A sky130_fd_sc_hd__and3_1
X_15973_ _15984_/CLK _15973_/D vssd1 vssd1 vccd1 vccd1 _15973_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10047_ _10047_/A _10047_/B vssd1 vssd1 vccd1 vccd1 _10048_/B sky130_fd_sc_hd__nor2_1
X_14924_ _14919_/A _14922_/B _14845_/X vssd1 vssd1 vccd1 vccd1 _14930_/C sky130_fd_sc_hd__o21a_1
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14855_ _14855_/A _14855_/B vssd1 vssd1 vccd1 vccd1 _16285_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13806_ _16070_/Q _13805_/C _13708_/X vssd1 vssd1 vccd1 vccd1 _13807_/B sky130_fd_sc_hd__a21oi_1
X_14786_ _14946_/A _14786_/B _14786_/C vssd1 vssd1 vccd1 vccd1 _14787_/A sky130_fd_sc_hd__and3_1
X_11998_ _11998_/A vssd1 vssd1 vccd1 vccd1 _15769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13737_ _14073_/A vssd1 vssd1 vccd1 vccd1 _13789_/A sky130_fd_sc_hd__clkbuf_2
X_10949_ _15607_/Q _10950_/B _10948_/X vssd1 vssd1 vccd1 vccd1 _10949_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15322_/CLK sky130_fd_sc_hd__clkbuf_16
X_13668_ _13666_/X _13664_/C _13667_/Y vssd1 vssd1 vccd1 vccd1 _16043_/D sky130_fd_sc_hd__a21oi_1
X_15407_ _15483_/CLK _15407_/D vssd1 vssd1 vccd1 vccd1 _15407_/Q sky130_fd_sc_hd__dfxtp_1
X_12619_ _12615_/X _12617_/Y _12618_/Y _12613_/C vssd1 vssd1 vccd1 vccd1 _12621_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13599_ _16033_/Q _13605_/C _13598_/X vssd1 vssd1 vccd1 vccd1 _13599_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15338_ _15339_/CLK _15338_/D vssd1 vssd1 vccd1 vccd1 _15338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_0 state1[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15269_ _15286_/CLK _15269_/D vssd1 vssd1 vccd1 vccd1 _15269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _13720_/A vssd1 vssd1 vccd1 vccd1 _10983_/A sky130_fd_sc_hd__clkbuf_4
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09761_ _09759_/A _09759_/B _09760_/X vssd1 vssd1 vccd1 vccd1 _15420_/D sky130_fd_sc_hd__a21oi_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08718_/A _08707_/Y _08711_/Y _08704_/C vssd1 vssd1 vccd1 vccd1 _08714_/B
+ sky130_fd_sc_hd__o211a_1
X_09692_ _15411_/Q _09867_/B _09692_/C vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__and3_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08643_ _15249_/Q _08872_/B _08651_/C vssd1 vssd1 vccd1 vccd1 _08643_/X sky130_fd_sc_hd__and3_1
XFILLER_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _10896_/A vssd1 vssd1 vccd1 vccd1 _13064_/B sky130_fd_sc_hd__buf_4
XFILLER_81_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16364_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ _15323_/Q _09125_/C _08888_/X vssd1 vssd1 vccd1 vccd1 _09127_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09057_ _09055_/Y _09050_/C _09052_/X _09053_/Y vssd1 vssd1 vccd1 vccd1 _09058_/C
+ sky130_fd_sc_hd__a211o_1
X_08008_ _13266_/C _13372_/C _08007_/Y vssd1 vssd1 vccd1 vccd1 _08010_/B sky130_fd_sc_hd__o21a_2
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09959_ _15453_/Q _09967_/C _09786_/X vssd1 vssd1 vccd1 vccd1 _09959_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_58_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12970_ _12977_/B _12970_/B vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__or2_1
XFILLER_58_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11921_ _11921_/A vssd1 vssd1 vccd1 vccd1 _15757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14640_ hold26/A _14639_/C _14095_/B vssd1 vssd1 vccd1 vccd1 _14641_/B sky130_fd_sc_hd__a21oi_1
X_11852_ _11885_/C vssd1 vssd1 vccd1 vccd1 _11891_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10803_ _10916_/A _10806_/C vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__or2_1
XFILLER_82_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14571_ _14565_/Y _14566_/X _14568_/B vssd1 vssd1 vccd1 vccd1 _14572_/B sky130_fd_sc_hd__o21a_1
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11783_ _11783_/A vssd1 vssd1 vccd1 vccd1 _12015_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_52_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16321_/CLK sky130_fd_sc_hd__clkbuf_16
X_16310_ _16317_/CLK _16310_/D vssd1 vssd1 vccd1 vccd1 _16310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13522_ _16020_/Q _13554_/C _13317_/X vssd1 vssd1 vccd1 vccd1 _13524_/B sky130_fd_sc_hd__a21oi_1
X_10734_ _15573_/Q _10734_/B _10734_/C vssd1 vssd1 vccd1 vccd1 _10744_/A sky130_fd_sc_hd__and3_1
XFILLER_15_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16241_ _16241_/CLK _16241_/D vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfxtp_1
X_13453_ _16007_/Q _13451_/C _13452_/X vssd1 vssd1 vccd1 vccd1 _13454_/B sky130_fd_sc_hd__a21oi_1
X_10665_ _15561_/Q _10778_/B _10665_/C vssd1 vssd1 vccd1 vccd1 _10665_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ _12518_/A _12404_/B _12408_/B vssd1 vssd1 vccd1 vccd1 _15833_/D sky130_fd_sc_hd__nor3_1
X_16172_ _16192_/CLK _16172_/D vssd1 vssd1 vccd1 vccd1 _16172_/Q sky130_fd_sc_hd__dfxtp_2
X_13384_ _13410_/A _13384_/B _13384_/C vssd1 vssd1 vccd1 vccd1 _13385_/A sky130_fd_sc_hd__and3_1
X_10596_ _15552_/Q _10654_/B _10596_/C vssd1 vssd1 vccd1 vccd1 _10596_/X sky130_fd_sc_hd__and3_1
XFILLER_139_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15123_ _14970_/X _15122_/A _15014_/X vssd1 vssd1 vccd1 vccd1 _15123_/Y sky130_fd_sc_hd__a21oi_1
X_12335_ _12331_/X _12333_/Y _12334_/Y _12329_/C vssd1 vssd1 vccd1 vccd1 _12337_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_5_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15054_ _14970_/X _15053_/A _15014_/X vssd1 vssd1 vccd1 vccd1 _15054_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12266_ _12281_/A _12266_/B _12266_/C vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__and3_1
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14005_ _16106_/Q _14003_/C _14004_/X vssd1 vssd1 vccd1 vccd1 _14006_/B sky130_fd_sc_hd__a21o_1
X_11217_ _15649_/Q _11259_/C _11047_/X vssd1 vssd1 vccd1 vccd1 _11220_/B sky130_fd_sc_hd__a21oi_1
X_12197_ _13041_/A vssd1 vssd1 vccd1 vccd1 _12197_/X sky130_fd_sc_hd__clkbuf_2
X_11148_ _11204_/A _11151_/C vssd1 vssd1 vccd1 vccd1 _11148_/X sky130_fd_sc_hd__or2_1
XFILLER_95_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11079_ _15627_/Q _11086_/C _10848_/X vssd1 vssd1 vccd1 vccd1 _11079_/Y sky130_fd_sc_hd__a21oi_1
X_15956_ _15956_/CLK _15956_/D vssd1 vssd1 vccd1 vccd1 _15956_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14907_ _14908_/B _14908_/C _14908_/A vssd1 vssd1 vccd1 vccd1 _14909_/B sky130_fd_sc_hd__a21o_1
X_15887_ _15907_/CLK _15887_/D vssd1 vssd1 vccd1 vccd1 _15887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14838_ _16286_/Q _14953_/B _14838_/C vssd1 vssd1 vccd1 vccd1 _14840_/A sky130_fd_sc_hd__and3_1
XFILLER_17_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14769_ _14853_/A _14811_/B _14769_/C vssd1 vssd1 vccd1 vccd1 _14771_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_43_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16192_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08290_ _08220_/A _08220_/B _08289_/X vssd1 vssd1 vccd1 vccd1 _08297_/A sky130_fd_sc_hd__a21bo_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09813_ _15428_/Q _09813_/B _09817_/C vssd1 vssd1 vccd1 vccd1 _09813_/Y sky130_fd_sc_hd__nand3_1
XFILLER_99_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09744_ _09740_/X _09742_/Y _09743_/Y _09738_/C vssd1 vssd1 vccd1 vccd1 _09746_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09675_ _09690_/A _09675_/B _09675_/C vssd1 vssd1 vccd1 vccd1 _09676_/A sky130_fd_sc_hd__and3_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08626_ _15247_/Q _08636_/C _08625_/X vssd1 vssd1 vccd1 vccd1 _08626_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08557_ _08557_/A _08557_/B _08557_/C vssd1 vssd1 vccd1 vccd1 _08558_/C sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_34_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16103_/CLK sky130_fd_sc_hd__clkbuf_16
X_08488_ _08488_/A _08488_/B _08488_/C vssd1 vssd1 vccd1 vccd1 _08489_/C sky130_fd_sc_hd__nand3_1
XFILLER_22_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10450_ _10456_/A _10447_/Y _10449_/Y _10444_/C vssd1 vssd1 vccd1 vccd1 _10452_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09109_ _09109_/A vssd1 vssd1 vccd1 vccd1 _15319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10381_ _15518_/Q _10609_/B _10389_/C vssd1 vssd1 vccd1 vccd1 _10381_/X sky130_fd_sc_hd__and3_1
XFILLER_109_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12120_ _12234_/A _12120_/B _12124_/B vssd1 vssd1 vccd1 vccd1 _15788_/D sky130_fd_sc_hd__nor3_1
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12051_ _12047_/X _12049_/Y _12050_/Y _12045_/C vssd1 vssd1 vccd1 vccd1 _12053_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11002_ _10996_/B _10997_/C _10999_/X _11000_/Y vssd1 vssd1 vccd1 vccd1 _11003_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15810_ _07603_/A _15810_/D vssd1 vssd1 vccd1 vccd1 _15810_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15741_ _15794_/CLK _15741_/D vssd1 vssd1 vccd1 vccd1 _15741_/Q sky130_fd_sc_hd__dfxtp_1
X_12953_ _12953_/A vssd1 vssd1 vccd1 vccd1 _15921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11904_ _11941_/A _11904_/B _11904_/C vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__and3_1
X_15672_ _15763_/CLK _15672_/D vssd1 vssd1 vccd1 vccd1 _15672_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12884_/A _12884_/B _12884_/C vssd1 vssd1 vccd1 vccd1 _12885_/C sky130_fd_sc_hd__nand3_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _16238_/Q _14639_/C _14503_/X vssd1 vssd1 vccd1 vccd1 _14626_/B sky130_fd_sc_hd__a21oi_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11835_ _11843_/B _11835_/B vssd1 vssd1 vccd1 vccd1 _11839_/A sky130_fd_sc_hd__or2_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _16129_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _16221_/Q _14593_/B _14554_/C vssd1 vssd1 vccd1 vccd1 _14561_/A sky130_fd_sc_hd__and3_1
XFILLER_13_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11766_ _11766_/A vssd1 vssd1 vccd1 vccd1 _15733_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13505_ _16016_/Q _13504_/C _13452_/X vssd1 vssd1 vccd1 vccd1 _13506_/B sky130_fd_sc_hd__a21oi_1
X_10717_ _10710_/B _10711_/C _10714_/X _10715_/Y vssd1 vssd1 vccd1 vccd1 _10718_/C
+ sky130_fd_sc_hd__a211o_1
X_14485_ _14482_/B _14481_/Y _14482_/A vssd1 vssd1 vccd1 vccd1 _14485_/Y sky130_fd_sc_hd__o21bai_1
X_11697_ _15723_/Q _11697_/B _11697_/C vssd1 vssd1 vccd1 vccd1 _11697_/Y sky130_fd_sc_hd__nand3_1
XFILLER_13_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16224_ _16224_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 _16224_/Q sky130_fd_sc_hd__dfxtp_1
X_13436_ _16005_/Q _13589_/B _13445_/C vssd1 vssd1 vccd1 vccd1 _13436_/X sky130_fd_sc_hd__and3_1
X_10648_ _11222_/A vssd1 vssd1 vccd1 vccd1 _10648_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16155_ _16166_/CLK _16155_/D vssd1 vssd1 vccd1 vccd1 _16155_/Q sky130_fd_sc_hd__dfxtp_2
X_13367_ _13868_/A vssd1 vssd1 vccd1 vccd1 _13476_/A sky130_fd_sc_hd__clkbuf_2
X_10579_ _10615_/A _10579_/B _10579_/C vssd1 vssd1 vccd1 vccd1 _10580_/A sky130_fd_sc_hd__and3_1
X_15106_ _15106_/A _15106_/B _15110_/B vssd1 vssd1 vccd1 vccd1 _16344_/D sky130_fd_sc_hd__nor3_1
XFILLER_114_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12318_ _15822_/Q _12326_/C _12093_/X vssd1 vssd1 vccd1 vccd1 _12318_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16086_ _16367_/CLK _16086_/D vssd1 vssd1 vccd1 vccd1 _16086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _15980_/Q _13297_/C _13194_/X vssd1 vssd1 vccd1 vccd1 _13299_/B sky130_fd_sc_hd__a21oi_1
XFILLER_142_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15037_ _16331_/Q _15036_/C _14917_/X vssd1 vssd1 vccd1 vccd1 _15038_/B sky130_fd_sc_hd__a21oi_1
X_12249_ _12249_/A vssd1 vssd1 vccd1 vccd1 _12262_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07790_ _15890_/Q vssd1 vssd1 vccd1 vccd1 _12763_/A sky130_fd_sc_hd__clkinv_2
XFILLER_84_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15939_ _15196_/Q _15939_/D vssd1 vssd1 vccd1 vccd1 _15939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09460_ _15375_/Q _09577_/B _09460_/C vssd1 vssd1 vccd1 vccd1 _09470_/A sky130_fd_sc_hd__and3_1
XFILLER_64_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ _08411_/A _08411_/B _08411_/C vssd1 vssd1 vccd1 vccd1 _08412_/C sky130_fd_sc_hd__or3_1
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09391_ _15363_/Q _09623_/B _09391_/C vssd1 vssd1 vccd1 vccd1 _09391_/Y sky130_fd_sc_hd__nand3_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _16040_/CLK sky130_fd_sc_hd__clkbuf_16
X_08342_ _08297_/A _08297_/B _08341_/X vssd1 vssd1 vccd1 vccd1 _08362_/A sky130_fd_sc_hd__a21bo_1
XFILLER_149_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08273_ _15209_/Q _08279_/A vssd1 vssd1 vccd1 vccd1 _08332_/B sky130_fd_sc_hd__and2_1
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07988_ _10347_/A _07827_/B _07826_/B vssd1 vssd1 vccd1 vccd1 _08042_/A sky130_fd_sc_hd__o21ai_2
XFILLER_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09727_ _15417_/Q _09784_/B _09727_/C vssd1 vssd1 vccd1 vccd1 _09727_/X sky130_fd_sc_hd__and3_1
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09658_ _09658_/A vssd1 vssd1 vccd1 vccd1 _09671_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _15245_/Q _08657_/C _07623_/X vssd1 vssd1 vccd1 vccd1 _08611_/B sky130_fd_sc_hd__a21oi_1
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09589_/A _09589_/B vssd1 vssd1 vccd1 vccd1 _09594_/C sky130_fd_sc_hd__nor2_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _15710_/Q vssd1 vssd1 vccd1 vccd1 _11635_/C sky130_fd_sc_hd__inv_2
XFILLER_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11551_ _11551_/A vssd1 vssd1 vccd1 vccd1 _11780_/A sky130_fd_sc_hd__clkbuf_2
X_10502_ _10500_/Y _10495_/C _10497_/X _10498_/Y vssd1 vssd1 vccd1 vccd1 _10503_/C
+ sky130_fd_sc_hd__a211o_1
X_14270_ _14270_/A vssd1 vssd1 vccd1 vccd1 _14270_/X sky130_fd_sc_hd__buf_2
X_11482_ _11491_/A _11480_/Y _11481_/Y _11477_/C vssd1 vssd1 vccd1 vccd1 _11484_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13221_ _13222_/B _13222_/C _13222_/A vssd1 vssd1 vccd1 vccd1 _13223_/B sky130_fd_sc_hd__a21o_1
X_10433_ _15526_/Q _10434_/C _10373_/X vssd1 vssd1 vccd1 vccd1 _10433_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13152_ _13617_/A vssd1 vssd1 vccd1 vccd1 _13666_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10364_ _10940_/A vssd1 vssd1 vccd1 vccd1 _10364_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _12099_/X _12101_/Y _12102_/Y _12097_/C vssd1 vssd1 vccd1 vccd1 _12105_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13199_/A _13086_/C vssd1 vssd1 vccd1 vccd1 _13083_/X sky130_fd_sc_hd__or2_1
X_10295_ _11507_/A vssd1 vssd1 vccd1 vccd1 _10532_/B sky130_fd_sc_hd__clkbuf_2
X_12034_ _15777_/Q _12042_/C _11805_/X vssd1 vssd1 vccd1 vccd1 _12034_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13985_ _13985_/A _13985_/B _13985_/C vssd1 vssd1 vccd1 vccd1 _13986_/C sky130_fd_sc_hd__nand3_1
X_15724_ _15794_/CLK _15724_/D vssd1 vssd1 vccd1 vccd1 _15724_/Q sky130_fd_sc_hd__dfxtp_1
X_12936_ _15920_/Q _12941_/C _13099_/A vssd1 vssd1 vccd1 vccd1 _12938_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15655_ _15655_/CLK _15655_/D vssd1 vssd1 vccd1 vccd1 _15655_/Q sky130_fd_sc_hd__dfxtp_1
X_12867_ _12865_/A _12865_/B _12866_/X vssd1 vssd1 vccd1 vccd1 _15906_/D sky130_fd_sc_hd__a21oi_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11818_ _11818_/A vssd1 vssd1 vccd1 vccd1 _15741_/D sky130_fd_sc_hd__clkbuf_1
X_14606_ _16232_/Q _14605_/C _07674_/A vssd1 vssd1 vccd1 vccd1 _14607_/B sky130_fd_sc_hd__a21o_1
X_15586_ _15194_/Q _15586_/D vssd1 vssd1 vccd1 vccd1 _15586_/Q sky130_fd_sc_hd__dfxtp_1
X_12798_ _15897_/Q _12798_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12808_/A sky130_fd_sc_hd__and3_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14537_ _07701_/X _14533_/B _14814_/A vssd1 vssd1 vccd1 vccd1 _14539_/A sky130_fd_sc_hd__a21oi_1
X_11749_ _11765_/A _11749_/B _11749_/C vssd1 vssd1 vccd1 vccd1 _11750_/A sky130_fd_sc_hd__and3_1
X_14468_ _16202_/Q _14468_/B _14474_/C vssd1 vssd1 vccd1 vccd1 _14471_/B sky130_fd_sc_hd__nand3_1
XFILLER_128_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13419_ _16002_/Q _13451_/C _13317_/X vssd1 vssd1 vccd1 vccd1 _13421_/B sky130_fd_sc_hd__a21oi_1
X_16207_ _16240_/CLK _16207_/D vssd1 vssd1 vccd1 vccd1 _16207_/Q sky130_fd_sc_hd__dfxtp_2
X_14399_ _14398_/X _14397_/Y _14309_/X vssd1 vssd1 vccd1 vccd1 _14399_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16138_ _16143_/CLK _16138_/D vssd1 vssd1 vccd1 vccd1 _16138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08960_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08999_/A sky130_fd_sc_hd__clkbuf_2
X_16069_ _16075_/CLK _16069_/D vssd1 vssd1 vccd1 vccd1 _16069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15961_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07911_ _15990_/Q vssd1 vssd1 vccd1 vccd1 _13420_/C sky130_fd_sc_hd__inv_4
X_08891_ _08891_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08892_/B sky130_fd_sc_hd__nor2_1
X_07842_ _07842_/A _07842_/B vssd1 vssd1 vccd1 vccd1 _07843_/B sky130_fd_sc_hd__nand2_2
XFILLER_111_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07773_ _16242_/Q vssd1 vssd1 vccd1 vccd1 _07777_/A sky130_fd_sc_hd__clkinv_2
X_09512_ _09512_/A vssd1 vssd1 vccd1 vccd1 _15381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _09443_/A vssd1 vssd1 vccd1 vccd1 _15371_/D sky130_fd_sc_hd__clkbuf_1
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09374_ _15362_/Q _09432_/B _09380_/C vssd1 vssd1 vccd1 vccd1 _09377_/B sky130_fd_sc_hd__nand3_1
X_08325_ _08325_/A _08339_/A vssd1 vssd1 vccd1 vccd1 _08326_/B sky130_fd_sc_hd__xor2_4
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08256_ _08256_/A _08256_/B vssd1 vssd1 vccd1 vccd1 _08256_/Y sky130_fd_sc_hd__nor2_1
X_08187_ _08187_/A _08187_/B vssd1 vssd1 vccd1 vccd1 _08191_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10080_ _10080_/A vssd1 vssd1 vccd1 vccd1 _15470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13770_ _13617_/X _13768_/C _13720_/X vssd1 vssd1 vccd1 vccd1 _13770_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10982_ _10982_/A vssd1 vssd1 vccd1 vccd1 _15610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12721_ _15885_/Q _12729_/C _12661_/X vssd1 vssd1 vccd1 vccd1 _12721_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ _15440_/CLK _15440_/D vssd1 vssd1 vccd1 vccd1 _15440_/Q sky130_fd_sc_hd__dfxtp_4
X_12652_ _12652_/A _12652_/B _12657_/A vssd1 vssd1 vccd1 vccd1 _15873_/D sky130_fd_sc_hd__nor3_1
XFILLER_130_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ _11601_/Y _11597_/C _11608_/A _11600_/Y vssd1 vssd1 vccd1 vccd1 _11608_/B
+ sky130_fd_sc_hd__a211oi_1
X_15371_ _15484_/CLK _15371_/D vssd1 vssd1 vccd1 vccd1 _15371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12583_ _12583_/A _12583_/B _12583_/C vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__or3_1
XFILLER_11_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14322_ _14190_/X _14320_/B _14321_/Y vssd1 vssd1 vccd1 vccd1 _16167_/D sky130_fd_sc_hd__o21a_1
X_11534_ _15698_/Q _11541_/C _11472_/X vssd1 vssd1 vccd1 vccd1 _11534_/Y sky130_fd_sc_hd__a21oi_1
X_14253_ _14253_/A _14253_/B _14253_/C vssd1 vssd1 vccd1 vccd1 _14254_/C sky130_fd_sc_hd__nand3_1
X_11465_ _12041_/A vssd1 vssd1 vccd1 vccd1 _11697_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_137_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _13223_/A _13204_/B _13204_/C vssd1 vssd1 vccd1 vccd1 _13205_/A sky130_fd_sc_hd__and3_1
X_10416_ _15523_/Q _10532_/B _10426_/C vssd1 vssd1 vccd1 vccd1 _10421_/A sky130_fd_sc_hd__and3_1
X_14184_ _14402_/A vssd1 vssd1 vccd1 vccd1 _14357_/B sky130_fd_sc_hd__clkbuf_2
X_11396_ _15677_/Q _11401_/C _11222_/X vssd1 vssd1 vccd1 vccd1 _11398_/C sky130_fd_sc_hd__a21o_1
X_13135_ _13133_/Y _13125_/C _13141_/A _13129_/Y vssd1 vssd1 vccd1 vccd1 _13141_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_124_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10347_ _10347_/A vssd1 vssd1 vccd1 vccd1 _10363_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _15941_/Q _13066_/B _13071_/C vssd1 vssd1 vccd1 vccd1 _13066_/Y sky130_fd_sc_hd__nand3_1
X_10278_ _10284_/B _10278_/B vssd1 vssd1 vccd1 vccd1 _10280_/A sky130_fd_sc_hd__or2_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12017_ _12053_/A _12017_/B _12017_/C vssd1 vssd1 vccd1 vccd1 _12018_/A sky130_fd_sc_hd__and3_1
XFILLER_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ _13925_/X _13964_/B _13926_/X vssd1 vssd1 vccd1 vccd1 _13971_/A sky130_fd_sc_hd__a21oi_1
XFILLER_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15707_ _15763_/CLK _15707_/D vssd1 vssd1 vccd1 vccd1 _15707_/Q sky130_fd_sc_hd__dfxtp_1
X_12919_ _12919_/A _12923_/C vssd1 vssd1 vccd1 vccd1 _12919_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13899_ _13896_/X _13895_/Y _14612_/A vssd1 vssd1 vccd1 vccd1 _13899_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15638_ _15728_/CLK _15638_/D vssd1 vssd1 vccd1 vccd1 _15638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _15655_/CLK _15569_/D vssd1 vssd1 vccd1 vccd1 _15569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _15096_/C _07735_/B _07739_/A vssd1 vssd1 vccd1 vccd1 _08115_/A sky130_fd_sc_hd__o21ai_4
XFILLER_30_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09090_ _15318_/Q _09146_/B _09096_/C vssd1 vssd1 vccd1 vccd1 _09093_/B sky130_fd_sc_hd__nand3_1
XFILLER_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08041_ _08041_/A _08041_/B vssd1 vssd1 vccd1 vccd1 _08042_/B sky130_fd_sc_hd__xor2_4
XFILLER_119_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09992_ _09992_/A _09992_/B vssd1 vssd1 vccd1 vccd1 _09993_/B sky130_fd_sc_hd__nor2_1
XFILLER_130_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ _08943_/A vssd1 vssd1 vccd1 vccd1 _15293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08874_ _15285_/Q _08880_/C _08873_/X vssd1 vssd1 vccd1 vccd1 _08874_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07825_ _15530_/Q _07825_/B vssd1 vssd1 vccd1 vccd1 _07826_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07756_ _13097_/C _07756_/B vssd1 vssd1 vccd1 vccd1 _07757_/B sky130_fd_sc_hd__xnor2_2
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07687_ _14806_/A vssd1 vssd1 vccd1 vccd1 _14964_/A sky130_fd_sc_hd__clkbuf_2
X_09426_ _09446_/C vssd1 vssd1 vccd1 vccd1 _09460_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09357_ _09357_/A _09357_/B vssd1 vssd1 vccd1 vccd1 _09358_/B sky130_fd_sc_hd__nor2_1
X_08308_ _08344_/A _08344_/B vssd1 vssd1 vccd1 vccd1 _08311_/A sky130_fd_sc_hd__xor2_1
XFILLER_138_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09288_ _09288_/A _09288_/B _09288_/C vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__and3_1
X_08239_ _08239_/A _08306_/A vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__xnor2_4
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _11250_/A vssd1 vssd1 vccd1 vccd1 _15652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10201_ _10199_/Y _10195_/C _10197_/X _10198_/Y vssd1 vssd1 vccd1 vccd1 _10202_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_109_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11181_ _11189_/A _11181_/B _11181_/C vssd1 vssd1 vccd1 vccd1 _11182_/A sky130_fd_sc_hd__and3_1
XFILLER_134_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10132_ _10153_/A _10132_/B _10132_/C vssd1 vssd1 vccd1 vccd1 _10133_/A sky130_fd_sc_hd__and3_1
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10063_ _15469_/Q _10239_/B _10074_/C vssd1 vssd1 vccd1 vccd1 _10071_/A sky130_fd_sc_hd__and3_1
XFILLER_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14940_ _15023_/A _14940_/B _14945_/A vssd1 vssd1 vccd1 vccd1 _16306_/D sky130_fd_sc_hd__nor3_1
XFILLER_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14871_ _16294_/Q _14875_/C _14789_/X vssd1 vssd1 vccd1 vccd1 _14871_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13822_ _14287_/A vssd1 vssd1 vccd1 vccd1 _13822_/X sky130_fd_sc_hd__buf_2
XFILLER_18_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13753_ _16060_/Q _13758_/C _13598_/X vssd1 vssd1 vccd1 vccd1 _13753_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10965_ _15608_/Q _10970_/B _10965_/C vssd1 vssd1 vccd1 vccd1 _10965_/Y sky130_fd_sc_hd__nand3_1
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ _13723_/A vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__clkbuf_4
X_13684_ _13735_/A _13684_/B _13684_/C vssd1 vssd1 vccd1 vccd1 _13685_/A sky130_fd_sc_hd__and3_1
XFILLER_16_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10896_ _10896_/A vssd1 vssd1 vccd1 vccd1 _12048_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15423_ _15483_/CLK _15423_/D vssd1 vssd1 vccd1 vccd1 _15423_/Q sky130_fd_sc_hd__dfxtp_2
X_12635_ _12635_/A _12635_/B vssd1 vssd1 vccd1 vccd1 _12640_/C sky130_fd_sc_hd__nor2_1
XFILLER_12_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15354_ _15356_/CLK _15354_/D vssd1 vssd1 vccd1 vccd1 _15354_/Q sky130_fd_sc_hd__dfxtp_1
X_12566_ _12566_/A vssd1 vssd1 vccd1 vccd1 _15859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11517_ _11517_/A vssd1 vssd1 vccd1 vccd1 _15694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14305_ _16168_/Q _14440_/B _14313_/C vssd1 vssd1 vccd1 vccd1 _14308_/A sky130_fd_sc_hd__and3_1
X_15285_ _15286_/CLK _15285_/D vssd1 vssd1 vccd1 vccd1 _15285_/Q sky130_fd_sc_hd__dfxtp_1
X_12497_ _12497_/A vssd1 vssd1 vccd1 vccd1 _15848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14236_ _14190_/X _14234_/B _14235_/Y vssd1 vssd1 vccd1 vccd1 _16149_/D sky130_fd_sc_hd__o21a_1
X_11448_ _15685_/Q _11487_/C _11336_/X vssd1 vssd1 vccd1 vccd1 _11450_/B sky130_fd_sc_hd__a21oi_1
XFILLER_109_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14167_ _14168_/B _14168_/C _14168_/A vssd1 vssd1 vccd1 vccd1 _14169_/B sky130_fd_sc_hd__a21o_1
X_11379_ _11493_/A _11382_/C vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__or2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13118_ _15951_/Q _13127_/C _15176_/B vssd1 vssd1 vccd1 vccd1 _13118_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_112_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14098_/A _14098_/B _14102_/B vssd1 vssd1 vccd1 vccd1 _16121_/D sky130_fd_sc_hd__nor3_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13069_/A _13049_/B _13049_/C vssd1 vssd1 vccd1 vccd1 _13050_/A sky130_fd_sc_hd__and3_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07610_ input9/X vssd1 vssd1 vccd1 vccd1 _13250_/A sky130_fd_sc_hd__buf_6
XFILLER_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08590_ _13078_/B vssd1 vssd1 vccd1 vccd1 _08590_/X sky130_fd_sc_hd__buf_2
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09211_ _15337_/Q _09211_/B _09211_/C vssd1 vssd1 vccd1 vccd1 _09211_/X sky130_fd_sc_hd__and3_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09142_ _15326_/Q _09179_/C _09029_/X vssd1 vssd1 vccd1 vccd1 _09145_/B sky130_fd_sc_hd__a21oi_1
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09073_ _09071_/A _09071_/B _09072_/X vssd1 vssd1 vccd1 vccd1 _15313_/D sky130_fd_sc_hd__a21oi_1
XFILLER_147_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08024_ _07822_/A _07822_/B _07821_/A vssd1 vssd1 vccd1 vccd1 _08214_/B sky130_fd_sc_hd__o21ai_2
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09975_ _09972_/X _09973_/Y _09974_/Y _09970_/C vssd1 vssd1 vccd1 vccd1 _09977_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08926_ input4/X vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__buf_4
XFILLER_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08857_ _08878_/A _08857_/B _08857_/C vssd1 vssd1 vccd1 vccd1 _08858_/A sky130_fd_sc_hd__and3_1
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07808_ _07808_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _07822_/A sky130_fd_sc_hd__nand2_2
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08788_ _08944_/A vssd1 vssd1 vccd1 vccd1 _08909_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07739_ _07739_/A _07739_/B vssd1 vssd1 vccd1 vccd1 _07740_/B sky130_fd_sc_hd__nand2_4
XFILLER_26_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10750_ _10863_/A _10750_/B _10750_/C vssd1 vssd1 vccd1 vccd1 _10753_/B sky130_fd_sc_hd__or3_1
XFILLER_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09409_ _09487_/A _09409_/B _09414_/B vssd1 vssd1 vccd1 vccd1 _15365_/D sky130_fd_sc_hd__nor3_1
XFILLER_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ _15563_/Q _10681_/B _10685_/C vssd1 vssd1 vccd1 vccd1 _10681_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _12420_/A vssd1 vssd1 vccd1 vccd1 _12434_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12351_ _12351_/A _12351_/B vssd1 vssd1 vccd1 vccd1 _12356_/C sky130_fd_sc_hd__nor2_1
XFILLER_126_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11302_ _11302_/A vssd1 vssd1 vccd1 vccd1 _15660_/D sky130_fd_sc_hd__clkbuf_1
X_15070_ _15064_/B _15065_/C _15075_/A _15068_/Y vssd1 vssd1 vccd1 vccd1 _15075_/B
+ sky130_fd_sc_hd__a211oi_1
X_12282_ _12282_/A vssd1 vssd1 vccd1 vccd1 _15814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14021_ _16111_/Q _14046_/C _13822_/X vssd1 vssd1 vccd1 vccd1 _14023_/B sky130_fd_sc_hd__a21oi_1
X_11233_ _11225_/B _11226_/C _11228_/X _11231_/Y vssd1 vssd1 vccd1 vccd1 _11234_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11164_ _15641_/Q _11169_/C _10933_/X vssd1 vssd1 vccd1 vccd1 _11166_/C sky130_fd_sc_hd__a21o_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10115_ _10284_/A _10115_/B _10115_/C vssd1 vssd1 vccd1 vccd1 _10117_/B sky130_fd_sc_hd__or3_1
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11095_ _11094_/B _11094_/C _11038_/X vssd1 vssd1 vccd1 vccd1 _11096_/C sky130_fd_sc_hd__o21ai_1
XFILLER_110_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15972_ _15984_/CLK _15972_/D vssd1 vssd1 vccd1 vccd1 _15972_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_103_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10046_ _10053_/B _10046_/B vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__or2_1
X_14923_ _14921_/A _14921_/B _14922_/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__a21oi_1
XFILLER_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14854_ _14694_/X _14851_/A _14808_/X vssd1 vssd1 vccd1 vccd1 _14855_/B sky130_fd_sc_hd__o21ai_1
XFILLER_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13805_ _16070_/Q _13853_/B _13805_/C vssd1 vssd1 vccd1 vccd1 _13812_/B sky130_fd_sc_hd__and3_1
X_11997_ _11997_/A _11997_/B _11997_/C vssd1 vssd1 vccd1 vccd1 _11998_/A sky130_fd_sc_hd__and3_1
X_14785_ _14785_/A _14785_/B _14785_/C vssd1 vssd1 vccd1 vccd1 _14786_/C sky130_fd_sc_hd__nand3_1
XFILLER_44_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13736_ _13736_/A vssd1 vssd1 vccd1 vccd1 _16055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10948_ _12100_/A vssd1 vssd1 vccd1 vccd1 _10948_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10879_ _10879_/A _10879_/B _10879_/C vssd1 vssd1 vccd1 vccd1 _10880_/C sky130_fd_sc_hd__nand3_1
X_13667_ _13617_/X _13664_/C _13464_/X vssd1 vssd1 vccd1 vccd1 _13667_/Y sky130_fd_sc_hd__o21ai_1
X_15406_ _15483_/CLK _15406_/D vssd1 vssd1 vccd1 vccd1 _15406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12618_ _15868_/Q _12793_/B _12623_/C vssd1 vssd1 vccd1 vccd1 _12618_/Y sky130_fd_sc_hd__nand3_1
X_13598_ _13598_/A vssd1 vssd1 vccd1 vccd1 _13598_/X sky130_fd_sc_hd__clkbuf_2
X_15337_ _15337_/CLK _15337_/D vssd1 vssd1 vccd1 vccd1 _15337_/Q sky130_fd_sc_hd__dfxtp_1
X_12549_ _12543_/B _12544_/C _12546_/X _12547_/Y vssd1 vssd1 vccd1 vccd1 _12550_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_1 state1[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _15286_/CLK _15268_/D vssd1 vssd1 vccd1 vccd1 _15268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14219_ _14212_/B _14213_/C _14223_/A _14217_/Y vssd1 vssd1 vccd1 vccd1 _14223_/B
+ sky130_fd_sc_hd__a211oi_1
X_15199_ _16359_/CLK _15199_/D vssd1 vssd1 vccd1 vccd1 _15199_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _09760_/A _09764_/C vssd1 vssd1 vccd1 vccd1 _09760_/X sky130_fd_sc_hd__or2_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _15258_/Q _08947_/B _08715_/C vssd1 vssd1 vccd1 vccd1 _08711_/Y sky130_fd_sc_hd__nand3_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _09691_/A vssd1 vssd1 vccd1 vccd1 _15409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08642_ _09801_/A vssd1 vssd1 vccd1 vccd1 _08872_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _15240_/Q _11080_/A _08582_/C vssd1 vssd1 vccd1 vccd1 _08573_/X sky130_fd_sc_hd__and3_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09125_ _15323_/Q _09354_/B _09125_/C vssd1 vssd1 vccd1 vccd1 _09133_/B sky130_fd_sc_hd__and3_1
X_09056_ _09052_/X _09053_/Y _09055_/Y _09050_/C vssd1 vssd1 vccd1 vccd1 _09058_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_135_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08007_ _15999_/Q _08007_/B vssd1 vssd1 vccd1 vccd1 _08007_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09958_ _15453_/Q _10074_/B _09958_/C vssd1 vssd1 vccd1 vccd1 _09958_/X sky130_fd_sc_hd__and3_1
X_08909_ _08909_/A _08909_/B _08916_/A vssd1 vssd1 vccd1 vccd1 _15289_/D sky130_fd_sc_hd__nor3_1
XFILLER_57_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09889_ _15440_/Q vssd1 vssd1 vccd1 vccd1 _09903_/C sky130_fd_sc_hd__inv_2
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11920_ _11941_/A _11920_/B _11920_/C vssd1 vssd1 vccd1 vccd1 _11921_/A sky130_fd_sc_hd__and3_1
XFILLER_100_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11851_ _11872_/C vssd1 vssd1 vccd1 vccd1 _11885_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_26_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10802_ _10802_/A _10802_/B vssd1 vssd1 vccd1 vccd1 _10806_/C sky130_fd_sc_hd__nor2_1
XFILLER_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14570_ _14565_/Y _14568_/X _14569_/Y vssd1 vssd1 vccd1 vccd1 _16220_/D sky130_fd_sc_hd__o21a_1
X_11782_ _11842_/A vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10733_ _10733_/A vssd1 vssd1 vccd1 vccd1 _15571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13521_ _13548_/C vssd1 vssd1 vccd1 vccd1 _13554_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16240_ _16240_/CLK _16240_/D vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
X_13452_ _14099_/B vssd1 vssd1 vccd1 vccd1 _13452_/X sky130_fd_sc_hd__buf_2
X_10664_ _15562_/Q _10665_/C _10663_/X vssd1 vssd1 vccd1 vccd1 _10664_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12403_ _12401_/Y _12396_/C _12408_/A _12400_/Y vssd1 vssd1 vccd1 vccd1 _12408_/B
+ sky130_fd_sc_hd__a211oi_1
X_16171_ _16192_/CLK _16171_/D vssd1 vssd1 vccd1 vccd1 _16171_/Q sky130_fd_sc_hd__dfxtp_2
X_13383_ _13377_/B _13378_/C _13380_/X _13381_/Y vssd1 vssd1 vccd1 vccd1 _13384_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ _10595_/A vssd1 vssd1 vccd1 vccd1 _15550_/D sky130_fd_sc_hd__clkbuf_1
X_12334_ _15823_/Q _12507_/B _12339_/C vssd1 vssd1 vccd1 vccd1 _12334_/Y sky130_fd_sc_hd__nand3_1
X_15122_ _15122_/A _15122_/B vssd1 vssd1 vccd1 vccd1 _16348_/D sky130_fd_sc_hd__nor2_1
XFILLER_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15053_ _15053_/A _15053_/B vssd1 vssd1 vccd1 vccd1 _16330_/D sky130_fd_sc_hd__nor2_1
X_12265_ _12259_/B _12260_/C _12262_/X _12263_/Y vssd1 vssd1 vccd1 vccd1 _12266_/C
+ sky130_fd_sc_hd__a211o_1
X_14004_ _14270_/A vssd1 vssd1 vccd1 vccd1 _14004_/X sky130_fd_sc_hd__clkbuf_2
X_11216_ _11253_/C vssd1 vssd1 vccd1 vccd1 _11259_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12196_ _12228_/C vssd1 vssd1 vccd1 vccd1 _12235_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_96_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ _11147_/A _11147_/B vssd1 vssd1 vccd1 vccd1 _11151_/C sky130_fd_sc_hd__nor2_1
XFILLER_68_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11078_ _15627_/Q _11078_/B _11078_/C vssd1 vssd1 vccd1 vccd1 _11089_/A sky130_fd_sc_hd__and3_1
X_15955_ _15956_/CLK _15955_/D vssd1 vssd1 vccd1 vccd1 _15955_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10029_ _15464_/Q _10029_/B _10037_/C vssd1 vssd1 vccd1 vccd1 _10029_/X sky130_fd_sc_hd__and3_1
XFILLER_76_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14906_ hold19/A _14905_/C _14744_/X vssd1 vssd1 vccd1 vccd1 _14908_/C sky130_fd_sc_hd__a21o_1
X_15886_ _15907_/CLK _15886_/D vssd1 vssd1 vccd1 vccd1 _15886_/Q sky130_fd_sc_hd__dfxtp_1
X_14837_ _14915_/A _14837_/B _14841_/B vssd1 vssd1 vccd1 vccd1 _16281_/D sky130_fd_sc_hd__nor3_1
XFILLER_91_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14768_ _14768_/A _14768_/B vssd1 vssd1 vccd1 vccd1 _16266_/D sky130_fd_sc_hd__nor2_1
XFILLER_16_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13719_ _13719_/A vssd1 vssd1 vccd1 vccd1 _16051_/D sky130_fd_sc_hd__clkbuf_1
X_14699_ _07707_/X _14697_/A _14698_/Y vssd1 vssd1 vccd1 vccd1 _16250_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09812_ _15429_/Q _09817_/C _09693_/X vssd1 vssd1 vccd1 vccd1 _09812_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ _15418_/Q _09862_/B _09748_/C vssd1 vssd1 vccd1 vccd1 _09743_/Y sky130_fd_sc_hd__nand3_1
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09674_ _09668_/B _09669_/C _09671_/X _09672_/Y vssd1 vssd1 vccd1 vccd1 _09675_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _13051_/B vssd1 vssd1 vccd1 vccd1 _08625_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08557_/B _08557_/C _08557_/A vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__a21o_1
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08487_ _08488_/B _08488_/C _08488_/A vssd1 vssd1 vccd1 vccd1 _08489_/B sky130_fd_sc_hd__a21o_1
XFILLER_11_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09108_ _09115_/A _09108_/B _09108_/C vssd1 vssd1 vccd1 vccd1 _09109_/A sky130_fd_sc_hd__and3_1
X_10380_ _11303_/A vssd1 vssd1 vccd1 vccd1 _10609_/B sky130_fd_sc_hd__clkbuf_2
X_09039_ _15310_/Q _09211_/B _09039_/C vssd1 vssd1 vccd1 vccd1 _09039_/X sky130_fd_sc_hd__and3_1
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ _15778_/Q _12223_/B _12055_/C vssd1 vssd1 vccd1 vccd1 _12050_/Y sky130_fd_sc_hd__nand3_1
XFILLER_104_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11001_ _10999_/X _11000_/Y _10996_/B _10997_/C vssd1 vssd1 vccd1 vccd1 _11003_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_89_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15740_ _15794_/CLK _15740_/D vssd1 vssd1 vccd1 vccd1 _15740_/Q sky130_fd_sc_hd__dfxtp_1
X_12952_ _12959_/A _12952_/B _12952_/C vssd1 vssd1 vccd1 vccd1 _12953_/A sky130_fd_sc_hd__and3_1
XFILLER_46_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11903_ _11901_/B _11901_/C _11902_/X vssd1 vssd1 vccd1 vccd1 _11904_/C sky130_fd_sc_hd__o21ai_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _15763_/CLK _15671_/D vssd1 vssd1 vccd1 vccd1 _15671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12884_/B _12884_/C _12884_/A vssd1 vssd1 vccd1 vccd1 _12885_/B sky130_fd_sc_hd__a21o_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14627_/C vssd1 vssd1 vccd1 vccd1 _14639_/C sky130_fd_sc_hd__clkbuf_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11834_ _15745_/Q _11833_/C _11775_/X vssd1 vssd1 vccd1 vccd1 _11835_/B sky130_fd_sc_hd__a21oi_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11765_ _11765_/A _11765_/B _11765_/C vssd1 vssd1 vccd1 vccd1 _11766_/A sky130_fd_sc_hd__and3_1
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14553_ _14553_/A vssd1 vssd1 vccd1 vccd1 _16217_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _10714_/X _10715_/Y _10710_/B _10711_/C vssd1 vssd1 vccd1 vccd1 _10718_/B
+ sky130_fd_sc_hd__o211ai_1
X_13504_ _16016_/Q _13605_/B _13504_/C vssd1 vssd1 vccd1 vccd1 _13512_/B sky130_fd_sc_hd__and3_1
XFILLER_147_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11696_ _15724_/Q _11697_/C _11526_/X vssd1 vssd1 vccd1 vccd1 _11696_/Y sky130_fd_sc_hd__a21oi_1
X_14484_ _14482_/A _14482_/B _14481_/Y _14483_/Y vssd1 vssd1 vccd1 vccd1 _16201_/D
+ sky130_fd_sc_hd__o31a_1
X_16223_ _16362_/CLK _16223_/D vssd1 vssd1 vccd1 vccd1 _16223_/Q sky130_fd_sc_hd__dfxtp_1
X_10647_ _15560_/Q _10876_/B _10654_/C vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__nand3_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ _13435_/A vssd1 vssd1 vccd1 vccd1 _16002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16154_ _16166_/CLK _16154_/D vssd1 vssd1 vccd1 vccd1 _16154_/Q sky130_fd_sc_hd__dfxtp_2
X_13366_ _14541_/A vssd1 vssd1 vccd1 vccd1 _13868_/A sky130_fd_sc_hd__clkbuf_4
X_10578_ _10577_/B _10577_/C _10464_/X vssd1 vssd1 vccd1 vccd1 _10579_/C sky130_fd_sc_hd__o21ai_1
XFILLER_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15105_ _15099_/B _15100_/C _15110_/A _15103_/Y vssd1 vssd1 vccd1 vccd1 _15110_/B
+ sky130_fd_sc_hd__a211oi_1
X_12317_ _15822_/Q _12434_/B _12317_/C vssd1 vssd1 vccd1 vccd1 _12317_/X sky130_fd_sc_hd__and3_1
X_16085_ _16367_/CLK _16085_/D vssd1 vssd1 vccd1 vccd1 _16085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13297_ _15980_/Q _13349_/B _13297_/C vssd1 vssd1 vccd1 vccd1 _13304_/B sky130_fd_sc_hd__and3_1
X_15036_ _16331_/Q _15142_/B _15036_/C vssd1 vssd1 vccd1 vccd1 _15038_/A sky130_fd_sc_hd__and3_1
X_12248_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12179_ _15799_/Q _12178_/C _12063_/X vssd1 vssd1 vccd1 vccd1 _12180_/B sky130_fd_sc_hd__a21oi_1
XFILLER_122_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15938_ _15196_/Q _15938_/D vssd1 vssd1 vccd1 vccd1 _15938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15869_ _15907_/CLK _15869_/D vssd1 vssd1 vccd1 vccd1 _15869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08410_ _08411_/A _08411_/C _08411_/B vssd1 vssd1 vccd1 vccd1 _08412_/B sky130_fd_sc_hd__o21ai_1
X_09390_ _10548_/A vssd1 vssd1 vccd1 vccd1 _09623_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08341_ _08341_/A _08298_/A vssd1 vssd1 vccd1 vccd1 _08341_/X sky130_fd_sc_hd__or2b_1
XFILLER_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08272_ _08272_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _08436_/A sky130_fd_sc_hd__xor2_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07987_ _10234_/A _07849_/B _07986_/X vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__o21ai_4
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09726_ _09726_/A vssd1 vssd1 vccd1 vccd1 _15415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09657_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__buf_2
XFILLER_83_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _08651_/C vssd1 vssd1 vccd1 vccd1 _08657_/C sky130_fd_sc_hd__clkbuf_2
X_09588_ _09588_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09589_/B sky130_fd_sc_hd__nor2_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _13972_/A vssd1 vssd1 vccd1 vccd1 _08580_/A sky130_fd_sc_hd__clkbuf_2
X_11550_ _11550_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _11552_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10501_ _10497_/X _10498_/Y _10500_/Y _10495_/C vssd1 vssd1 vccd1 vccd1 _10503_/B
+ sky130_fd_sc_hd__o211ai_1
X_11481_ _15689_/Q _11601_/B _11487_/C vssd1 vssd1 vccd1 vccd1 _11481_/Y sky130_fd_sc_hd__nand3_1
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13220_ _15967_/Q _13226_/C _14250_/A vssd1 vssd1 vccd1 vccd1 _13222_/C sky130_fd_sc_hd__a21o_1
X_10432_ _15526_/Q _10602_/B _10434_/C vssd1 vssd1 vccd1 vccd1 _10432_/X sky130_fd_sc_hd__and3_1
XFILLER_109_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13151_ _13151_/A vssd1 vssd1 vccd1 vccd1 _13617_/A sky130_fd_sc_hd__clkinv_2
XFILLER_109_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ _15516_/Q _10363_/B _10363_/C vssd1 vssd1 vccd1 vccd1 _10363_/X sky130_fd_sc_hd__and3_1
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12102_ _15786_/Q _12270_/B _12102_/C vssd1 vssd1 vccd1 vccd1 _12102_/Y sky130_fd_sc_hd__nand3_1
X_13082_ _13082_/A _13082_/B vssd1 vssd1 vccd1 vccd1 _13086_/C sky130_fd_sc_hd__nor2_1
X_10294_ input1/X vssd1 vssd1 vccd1 vccd1 _11507_/A sky130_fd_sc_hd__buf_2
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12033_ _15777_/Q _12150_/B _12033_/C vssd1 vssd1 vccd1 vccd1 _12033_/X sky130_fd_sc_hd__and3_1
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13984_ _13985_/B _13985_/C _13985_/A vssd1 vssd1 vccd1 vccd1 _13986_/B sky130_fd_sc_hd__a21o_1
XFILLER_19_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15723_ _15794_/CLK _15723_/D vssd1 vssd1 vccd1 vccd1 _15723_/Q sky130_fd_sc_hd__dfxtp_1
X_12935_ _15920_/Q _12935_/B _12941_/C vssd1 vssd1 vccd1 vccd1 _12938_/B sky130_fd_sc_hd__nand3_1
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15654_ _15655_/CLK _15654_/D vssd1 vssd1 vccd1 vccd1 _15654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12866_ _12919_/A _12869_/C vssd1 vssd1 vccd1 vccd1 _12866_/X sky130_fd_sc_hd__or2_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _16232_/Q _14605_/B _14605_/C vssd1 vssd1 vccd1 vccd1 _14605_/X sky130_fd_sc_hd__and3_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11817_ _11824_/A _11817_/B _11817_/C vssd1 vssd1 vccd1 vccd1 _11818_/A sky130_fd_sc_hd__and3_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _15194_/Q _15585_/D vssd1 vssd1 vccd1 vccd1 _15585_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12797_/A vssd1 vssd1 vccd1 vccd1 _15895_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _14413_/X _14533_/B _14535_/Y vssd1 vssd1 vccd1 vccd1 _16213_/D sky130_fd_sc_hd__o21a_1
X_11748_ _11742_/B _11743_/C _11745_/X _11746_/Y vssd1 vssd1 vccd1 vccd1 _11749_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_146_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14467_ _14517_/A _14467_/B _14471_/A vssd1 vssd1 vccd1 vccd1 _16198_/D sky130_fd_sc_hd__nor3_1
X_11679_ _11712_/C vssd1 vssd1 vccd1 vccd1 _11719_/C sky130_fd_sc_hd__clkbuf_2
X_16206_ _16362_/CLK _16206_/D vssd1 vssd1 vccd1 vccd1 _16206_/Q sky130_fd_sc_hd__dfxtp_1
X_13418_ _13445_/C vssd1 vssd1 vccd1 vccd1 _13451_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14398_ _14398_/A _14398_/B vssd1 vssd1 vccd1 vccd1 _14398_/X sky130_fd_sc_hd__or2_1
X_16137_ _16148_/CLK _16137_/D vssd1 vssd1 vccd1 vccd1 _16137_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13349_ _15989_/Q _13349_/B _13349_/C vssd1 vssd1 vccd1 vccd1 _13358_/B sky130_fd_sc_hd__and3_1
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16068_ _16075_/CLK _16068_/D vssd1 vssd1 vccd1 vccd1 _16068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07910_ _15764_/Q _07957_/B vssd1 vssd1 vccd1 vccd1 _07920_/A sky130_fd_sc_hd__xnor2_4
X_15019_ _15024_/C vssd1 vssd1 vccd1 vccd1 _15036_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08890_ _08897_/B _08890_/B vssd1 vssd1 vccd1 vccd1 _08892_/A sky130_fd_sc_hd__or2_1
XFILLER_111_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07841_ _15917_/Q _15935_/Q vssd1 vssd1 vccd1 vccd1 _07842_/B sky130_fd_sc_hd__or2_1
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07772_ _07772_/A _08069_/B vssd1 vssd1 vccd1 vccd1 _07780_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ _09519_/A _09511_/B _09511_/C vssd1 vssd1 vccd1 vccd1 _09512_/A sky130_fd_sc_hd__and3_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09442_ _09458_/A _09442_/B _09442_/C vssd1 vssd1 vccd1 vccd1 _09443_/A sky130_fd_sc_hd__and3_1
XFILLER_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _09487_/A _09373_/B _09377_/A vssd1 vssd1 vccd1 vccd1 _15360_/D sky130_fd_sc_hd__nor3_1
XFILLER_33_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08324_ _08324_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08339_/A sky130_fd_sc_hd__xnor2_2
X_08255_ _08255_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__xnor2_4
XFILLER_119_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08186_ _08021_/A _08021_/B _08020_/A vssd1 vssd1 vccd1 vccd1 _08193_/A sky130_fd_sc_hd__a21o_2
XFILLER_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ _09708_/B _09708_/C _09596_/X vssd1 vssd1 vccd1 vccd1 _09710_/C sky130_fd_sc_hd__o21ai_1
XFILLER_74_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10981_ _11019_/A _10981_/B _10981_/C vssd1 vssd1 vccd1 vccd1 _10982_/A sky130_fd_sc_hd__and3_1
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12720_ _15885_/Q _12720_/B _12720_/C vssd1 vssd1 vccd1 vccd1 _12720_/X sky130_fd_sc_hd__and3_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12651_ _15874_/Q _12879_/B _12660_/C vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__and3_1
X_11602_ _11608_/A _11600_/Y _11601_/Y _11597_/C vssd1 vssd1 vccd1 vccd1 _11604_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15370_ _15484_/CLK _15370_/D vssd1 vssd1 vccd1 vccd1 _15370_/Q sky130_fd_sc_hd__dfxtp_1
X_12582_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12621_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14321_ _14321_/A _14321_/B vssd1 vssd1 vccd1 vccd1 _14321_/Y sky130_fd_sc_hd__nor2_1
X_11533_ _15698_/Q _11533_/B _11541_/C vssd1 vssd1 vccd1 vccd1 _11533_/X sky130_fd_sc_hd__and3_1
XFILLER_128_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14252_ _14253_/B _14253_/C _14253_/A vssd1 vssd1 vccd1 vccd1 _14254_/B sky130_fd_sc_hd__a21o_1
X_11464_ _15688_/Q _11466_/C _11237_/X vssd1 vssd1 vccd1 vccd1 _11464_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _15523_/Q _10453_/C _10181_/X vssd1 vssd1 vccd1 vccd1 _10417_/B sky130_fd_sc_hd__a21oi_1
X_13203_ _13202_/B _13202_/C _14892_/A vssd1 vssd1 vccd1 vccd1 _13204_/C sky130_fd_sc_hd__o21ai_1
XFILLER_137_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11395_ _15677_/Q _11510_/B _11401_/C vssd1 vssd1 vccd1 vccd1 _11398_/B sky130_fd_sc_hd__nand3_1
X_14183_ _14180_/B _14179_/Y _14180_/A vssd1 vssd1 vccd1 vccd1 _14183_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_125_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10346_ _15520_/Q _15519_/Q _15518_/Q _10119_/X vssd1 vssd1 vccd1 vccd1 _15512_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13134_ _13141_/A _13129_/Y _13133_/Y _13125_/C vssd1 vssd1 vccd1 vccd1 _13136_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13065_ _15942_/Q _13071_/C _07672_/A vssd1 vssd1 vccd1 vccd1 _13065_/Y sky130_fd_sc_hd__a21oi_1
X_10277_ _15502_/Q _10276_/C _10044_/X vssd1 vssd1 vccd1 vccd1 _10278_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12016_ _12015_/B _12015_/C _11902_/X vssd1 vssd1 vccd1 vccd1 _12017_/C sky130_fd_sc_hd__o21ai_1
XFILLER_39_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13967_ _13920_/X _13964_/B _13966_/Y vssd1 vssd1 vccd1 vccd1 _16096_/D sky130_fd_sc_hd__o21a_1
XFILLER_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15706_ _15794_/CLK _15706_/D vssd1 vssd1 vccd1 vccd1 _15706_/Q sky130_fd_sc_hd__dfxtp_1
X_12918_ _12918_/A _12918_/B vssd1 vssd1 vccd1 vccd1 _12923_/C sky130_fd_sc_hd__nor2_1
XFILLER_62_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13898_ _14883_/A vssd1 vssd1 vccd1 vccd1 _14612_/A sky130_fd_sc_hd__buf_2
XFILLER_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15637_ _15194_/Q _15637_/D vssd1 vssd1 vccd1 vccd1 _15637_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12849_ _12845_/X _12846_/Y _12848_/Y _12843_/C vssd1 vssd1 vccd1 vccd1 _12851_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15568_ _15655_/CLK _15568_/D vssd1 vssd1 vccd1 vccd1 _15568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14519_ _16213_/Q _14525_/C _14395_/X vssd1 vssd1 vccd1 vccd1 _14521_/B sky130_fd_sc_hd__a21oi_1
X_15499_ _15224_/Q _15499_/D vssd1 vssd1 vccd1 vccd1 _15499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08041_/B sky130_fd_sc_hd__xor2_4
XFILLER_134_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ _09997_/B _09991_/B vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__or2_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08942_ _08942_/A _08942_/B _08942_/C vssd1 vssd1 vccd1 vccd1 _08943_/A sky130_fd_sc_hd__and3_1
XFILLER_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08873_ _13064_/B vssd1 vssd1 vccd1 vccd1 _08873_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07824_ _15530_/Q _07825_/B vssd1 vssd1 vccd1 vccd1 _07826_/A sky130_fd_sc_hd__or2_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07755_ _07755_/A _07755_/B vssd1 vssd1 vccd1 vccd1 _07756_/B sky130_fd_sc_hd__nand2_2
XFILLER_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07686_ _14765_/A _07698_/C vssd1 vssd1 vccd1 vccd1 _07692_/A sky130_fd_sc_hd__and2_1
XFILLER_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ _09438_/C vssd1 vssd1 vccd1 vccd1 _09446_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09356_ _09362_/B _09356_/B vssd1 vssd1 vccd1 vccd1 _09358_/A sky130_fd_sc_hd__or2_1
XFILLER_100_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ _08238_/A _08238_/B _08306_/X vssd1 vssd1 vccd1 vccd1 _08344_/B sky130_fd_sc_hd__o21a_1
X_09287_ _09285_/Y _09281_/C _09283_/X _09284_/Y vssd1 vssd1 vccd1 vccd1 _09288_/C
+ sky130_fd_sc_hd__a211o_1
X_08238_ _08238_/A _08238_/B vssd1 vssd1 vccd1 vccd1 _08306_/A sky130_fd_sc_hd__xnor2_2
XFILLER_20_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08169_ _07946_/C _08166_/Y _08168_/X vssd1 vssd1 vccd1 vccd1 _08169_/Y sky130_fd_sc_hd__a21oi_1
X_10200_ _10197_/X _10198_/Y _10199_/Y _10195_/C vssd1 vssd1 vccd1 vccd1 _10202_/B
+ sky130_fd_sc_hd__o211ai_1
X_11180_ _11178_/Y _11173_/C _11175_/X _11176_/Y vssd1 vssd1 vccd1 vccd1 _11181_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10131_ _10131_/A _10131_/B _10131_/C vssd1 vssd1 vccd1 vccd1 _10132_/C sky130_fd_sc_hd__nand3_1
XFILLER_133_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10062_ _15469_/Q _10106_/C _09893_/X vssd1 vssd1 vccd1 vccd1 _10064_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14870_ _16294_/Q _15031_/B _14875_/C vssd1 vssd1 vccd1 vccd1 _14878_/A sky130_fd_sc_hd__and3_1
XFILLER_85_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13821_ _13846_/C vssd1 vssd1 vccd1 vccd1 _13853_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13752_ _16060_/Q _14093_/B _13752_/C vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__and3_1
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10964_ _15609_/Q _10970_/B _10848_/X vssd1 vssd1 vccd1 vccd1 _10964_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12703_ _13720_/A vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__buf_2
X_13683_ _13683_/A _13683_/B _13683_/C vssd1 vssd1 vccd1 vccd1 _13684_/C sky130_fd_sc_hd__nand3_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10895_ _15599_/Q _10895_/B _10904_/C vssd1 vssd1 vccd1 vccd1 _10895_/X sky130_fd_sc_hd__and3_1
X_15422_ _15422_/CLK _15422_/D vssd1 vssd1 vccd1 vccd1 _15422_/Q sky130_fd_sc_hd__dfxtp_2
X_12634_ _12634_/A _12634_/B vssd1 vssd1 vccd1 vccd1 _12635_/B sky130_fd_sc_hd__nor2_1
XFILLER_129_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15353_ _15356_/CLK _15353_/D vssd1 vssd1 vccd1 vccd1 _15353_/Q sky130_fd_sc_hd__dfxtp_1
X_12565_ _12565_/A _12565_/B _12565_/C vssd1 vssd1 vccd1 vccd1 _12566_/A sky130_fd_sc_hd__and3_1
XFILLER_129_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14304_ _14304_/A _14304_/B _14307_/B vssd1 vssd1 vccd1 vccd1 _16164_/D sky130_fd_sc_hd__nor3_1
X_11516_ _11538_/A _11516_/B _11516_/C vssd1 vssd1 vccd1 vccd1 _11517_/A sky130_fd_sc_hd__and3_1
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15284_ _15286_/CLK _15284_/D vssd1 vssd1 vccd1 vccd1 _15284_/Q sky130_fd_sc_hd__dfxtp_1
X_12496_ _12510_/A _12496_/B _12496_/C vssd1 vssd1 vccd1 vccd1 _12497_/A sky130_fd_sc_hd__and3_1
X_14235_ _14321_/A _14235_/B vssd1 vssd1 vccd1 vccd1 _14235_/Y sky130_fd_sc_hd__nor2_1
X_11447_ _11479_/C vssd1 vssd1 vccd1 vccd1 _11487_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11378_ _11378_/A _11378_/B vssd1 vssd1 vccd1 vccd1 _11382_/C sky130_fd_sc_hd__nor2_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14166_ _16139_/Q _14171_/C _13982_/X vssd1 vssd1 vccd1 vccd1 _14168_/C sky130_fd_sc_hd__a21o_1
XFILLER_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10329_ _10327_/Y _10323_/C _10336_/A _10326_/Y vssd1 vssd1 vccd1 vccd1 _10336_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _15951_/Q _13333_/B _13127_/C vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__and3_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14097_ _14095_/Y _14091_/C _14102_/A _14094_/Y vssd1 vssd1 vccd1 vccd1 _14102_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _13048_/A _13048_/B _13048_/C vssd1 vssd1 vccd1 vccd1 _13049_/C sky130_fd_sc_hd__nand3_1
XFILLER_112_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14999_ _15041_/A _14999_/B vssd1 vssd1 vccd1 vccd1 _14999_/X sky130_fd_sc_hd__or2_1
XFILLER_35_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09210_ _09210_/A vssd1 vssd1 vccd1 vccd1 _15335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09141_ _09173_/C vssd1 vssd1 vccd1 vccd1 _09179_/C sky130_fd_sc_hd__clkbuf_2
X_09072_ _09185_/A _09075_/C vssd1 vssd1 vccd1 vccd1 _09072_/X sky130_fd_sc_hd__or2_1
X_08023_ _12420_/A _07846_/B _08022_/Y vssd1 vssd1 vccd1 vccd1 _08037_/A sky130_fd_sc_hd__o21ai_4
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _15454_/Q _10150_/B _09979_/C vssd1 vssd1 vccd1 vccd1 _09974_/Y sky130_fd_sc_hd__nand3_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08925_ _08925_/A vssd1 vssd1 vccd1 vccd1 _15291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08856_ _08856_/A _08856_/B _08856_/C vssd1 vssd1 vccd1 vccd1 _08857_/C sky130_fd_sc_hd__nand3_1
X_07807_ _14289_/C _07807_/B vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__or2_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08787_ _15287_/Q _15286_/Q _15285_/Q _08604_/X vssd1 vssd1 vccd1 vccd1 _15270_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07738_ _15024_/C _07738_/B vssd1 vssd1 vccd1 vccd1 _07739_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07669_ _07667_/A _07667_/B _07668_/X vssd1 vssd1 vccd1 vccd1 _15201_/D sky130_fd_sc_hd__a21oi_1
XFILLER_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09408_ _09406_/Y _09401_/C _09414_/A _09405_/Y vssd1 vssd1 vccd1 vccd1 _09414_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_41_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10680_ _15564_/Q _10685_/C _10562_/X vssd1 vssd1 vccd1 vccd1 _10680_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09339_ _15357_/Q _09451_/B _09348_/C vssd1 vssd1 vccd1 vccd1 _09339_/X sky130_fd_sc_hd__and3_1
XFILLER_138_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12350_ _12350_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12351_/B sky130_fd_sc_hd__nor2_1
X_11301_ _11309_/A _11301_/B _11301_/C vssd1 vssd1 vccd1 vccd1 _11302_/A sky130_fd_sc_hd__and3_1
X_12281_ _12281_/A _12281_/B _12281_/C vssd1 vssd1 vccd1 vccd1 _12282_/A sky130_fd_sc_hd__and3_1
XFILLER_126_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _11228_/X _11231_/Y _11225_/B _11226_/C vssd1 vssd1 vccd1 vccd1 _11234_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_5_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14020_ _14032_/C vssd1 vssd1 vccd1 vccd1 _14046_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11163_ _15641_/Q _11221_/B _11169_/C vssd1 vssd1 vccd1 vccd1 _11166_/B sky130_fd_sc_hd__nand3_1
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10114_ _10114_/A vssd1 vssd1 vccd1 vccd1 _10153_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11094_ _11151_/A _11094_/B _11094_/C vssd1 vssd1 vccd1 vccd1 _11096_/B sky130_fd_sc_hd__or3_1
XFILLER_110_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15971_ _15971_/CLK _15971_/D vssd1 vssd1 vccd1 vccd1 _15971_/Q sky130_fd_sc_hd__dfxtp_1
X_10045_ _15466_/Q _10043_/C _10044_/X vssd1 vssd1 vccd1 vccd1 _10046_/B sky130_fd_sc_hd__a21oi_1
X_14922_ _15041_/A _14922_/B vssd1 vssd1 vccd1 vccd1 _14922_/X sky130_fd_sc_hd__or2_1
XFILLER_102_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14853_ _14853_/A _15010_/B _14853_/C vssd1 vssd1 vccd1 vccd1 _14855_/A sky130_fd_sc_hd__and3_1
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13804_ _13852_/A _13804_/B _13808_/B vssd1 vssd1 vccd1 vccd1 _16067_/D sky130_fd_sc_hd__nor3_1
XFILLER_16_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14784_ _14785_/B _14785_/C _14785_/A vssd1 vssd1 vccd1 vccd1 _14786_/B sky130_fd_sc_hd__a21o_1
X_11996_ _11994_/Y _11989_/C _11991_/X _11992_/Y vssd1 vssd1 vccd1 vccd1 _11997_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_91_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13735_ _13735_/A _13735_/B _13735_/C vssd1 vssd1 vccd1 vccd1 _13736_/A sky130_fd_sc_hd__and3_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10947_ _10947_/A vssd1 vssd1 vccd1 vccd1 _12100_/A sky130_fd_sc_hd__buf_6
X_13666_ _13666_/A vssd1 vssd1 vccd1 vccd1 _13666_/X sky130_fd_sc_hd__clkbuf_2
X_10878_ _10879_/B _10879_/C _10879_/A vssd1 vssd1 vccd1 vccd1 _10880_/B sky130_fd_sc_hd__a21o_1
X_15405_ _15483_/CLK _15405_/D vssd1 vssd1 vccd1 vccd1 _15405_/Q sky130_fd_sc_hd__dfxtp_2
X_12617_ _15869_/Q _12623_/C _12616_/X vssd1 vssd1 vccd1 vccd1 _12617_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13597_ _16033_/Q _13648_/B _13597_/C vssd1 vssd1 vccd1 vccd1 _13608_/A sky130_fd_sc_hd__and3_1
X_15336_ _15348_/CLK _15336_/D vssd1 vssd1 vccd1 vccd1 _15336_/Q sky130_fd_sc_hd__dfxtp_1
X_12548_ _12546_/X _12547_/Y _12543_/B _12544_/C vssd1 vssd1 vccd1 vccd1 _12550_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_129_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15267_ _15286_/CLK _15267_/D vssd1 vssd1 vccd1 vccd1 _15267_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_2 state1[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12500_/C vssd1 vssd1 vccd1 vccd1 _12512_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14218_ _14223_/A _14217_/Y _14212_/B _14213_/C vssd1 vssd1 vccd1 vccd1 _14220_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15198_ _16364_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 _15198_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14149_ _14368_/A vssd1 vssd1 vccd1 vccd1 _14149_/X sky130_fd_sc_hd__clkbuf_2
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _13598_/A vssd1 vssd1 vccd1 vccd1 _08947_/B sky130_fd_sc_hd__clkbuf_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _09690_/A _09690_/B _09690_/C vssd1 vssd1 vccd1 vccd1 _09691_/A sky130_fd_sc_hd__and3_1
XFILLER_67_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08641_ _10896_/A vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__buf_4
XFILLER_94_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08572_ _08572_/A vssd1 vssd1 vccd1 vccd1 _15238_/D sky130_fd_sc_hd__clkbuf_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09124_ _09699_/A vssd1 vssd1 vccd1 vccd1 _09354_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_148_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _15311_/Q _09285_/B _09061_/C vssd1 vssd1 vccd1 vccd1 _09055_/Y sky130_fd_sc_hd__nand3_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16370__19 vssd1 vssd1 vccd1 vccd1 _16370__19/HI io_oeb[2] sky130_fd_sc_hd__conb_1
X_08006_ _15981_/Q vssd1 vssd1 vccd1 vccd1 _13372_/C sky130_fd_sc_hd__inv_2
XFILLER_144_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_4_0_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_0_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_09957_ _09957_/A vssd1 vssd1 vccd1 vccd1 _15451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08908_ _15290_/Q _09088_/B _08919_/C vssd1 vssd1 vccd1 vccd1 _08916_/A sky130_fd_sc_hd__and3_1
X_09888_ _15448_/Q _15447_/Q _15446_/Q _09831_/X vssd1 vssd1 vccd1 vccd1 _15440_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08839_ _08839_/A _08839_/B _08839_/C vssd1 vssd1 vccd1 vccd1 _08841_/B sky130_fd_sc_hd__or3_1
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11850_ _11863_/C vssd1 vssd1 vccd1 vccd1 _11872_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10801_ _10801_/A _10801_/B vssd1 vssd1 vccd1 vccd1 _10802_/B sky130_fd_sc_hd__nor2_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11781_ _11779_/A _11779_/B _11780_/X vssd1 vssd1 vccd1 vccd1 _15735_/D sky130_fd_sc_hd__a21oi_1
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13520_ _13533_/C vssd1 vssd1 vccd1 vccd1 _13548_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10732_ _10732_/A _10732_/B _10732_/C vssd1 vssd1 vccd1 vccd1 _10733_/A sky130_fd_sc_hd__and3_1
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13451_ _16007_/Q _13605_/B _13451_/C vssd1 vssd1 vccd1 vccd1 _13460_/B sky130_fd_sc_hd__and3_1
X_10663_ _10663_/A vssd1 vssd1 vccd1 vccd1 _10663_/X sky130_fd_sc_hd__buf_2
X_12402_ _12408_/A _12400_/Y _12401_/Y _12396_/C vssd1 vssd1 vccd1 vccd1 _12404_/B
+ sky130_fd_sc_hd__o211a_1
X_16170_ _16204_/CLK _16170_/D vssd1 vssd1 vccd1 vccd1 _16170_/Q sky130_fd_sc_hd__dfxtp_1
X_10594_ _10615_/A _10594_/B _10594_/C vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__and3_1
X_13382_ _13380_/X _13381_/Y _13377_/B _13378_/C vssd1 vssd1 vccd1 vccd1 _13384_/B
+ sky130_fd_sc_hd__o211ai_1
X_15121_ _13920_/A _15119_/A _15086_/X vssd1 vssd1 vccd1 vccd1 _15122_/B sky130_fd_sc_hd__o21ai_1
X_12333_ _15824_/Q _12339_/C _12332_/X vssd1 vssd1 vccd1 vccd1 _12333_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_15052_ _14892_/X _15049_/A _15007_/X vssd1 vssd1 vccd1 vccd1 _15053_/B sky130_fd_sc_hd__o21ai_1
X_12264_ _12262_/X _12263_/Y _12259_/B _12260_/C vssd1 vssd1 vccd1 vccd1 _12266_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14003_ _16106_/Q _14137_/B _14003_/C vssd1 vssd1 vccd1 vccd1 _14003_/X sky130_fd_sc_hd__and3_1
X_11215_ _11239_/C vssd1 vssd1 vccd1 vccd1 _11253_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12195_ _12216_/C vssd1 vssd1 vccd1 vccd1 _12228_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11146_ _11146_/A _11146_/B vssd1 vssd1 vccd1 vccd1 _11147_/B sky130_fd_sc_hd__nor2_1
XFILLER_122_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11077_ _11077_/A vssd1 vssd1 vccd1 vccd1 _15625_/D sky130_fd_sc_hd__clkbuf_1
X_15954_ _15970_/CLK _15954_/D vssd1 vssd1 vccd1 vccd1 _15954_/Q sky130_fd_sc_hd__dfxtp_4
X_10028_ _10028_/A vssd1 vssd1 vccd1 vccd1 _15462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14905_ hold19/X _14941_/B _14905_/C vssd1 vssd1 vccd1 vccd1 _14908_/B sky130_fd_sc_hd__nand3_1
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15885_ _15907_/CLK _15885_/D vssd1 vssd1 vccd1 vccd1 _15885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14836_ _14829_/B _14830_/C _14841_/A _14834_/Y vssd1 vssd1 vccd1 vccd1 _14841_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14767_ _14766_/X _14769_/C _14695_/X vssd1 vssd1 vccd1 vccd1 _14768_/B sky130_fd_sc_hd__o21ai_1
X_11979_ _15768_/Q _11986_/C _11805_/X vssd1 vssd1 vccd1 vccd1 _11979_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13718_ _13735_/A _13718_/B _13718_/C vssd1 vssd1 vccd1 vccd1 _13719_/A sky130_fd_sc_hd__and3_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14698_ _07710_/X _14697_/A _14614_/X vssd1 vssd1 vccd1 vccd1 _14698_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13649_ _16042_/Q _13655_/C _13598_/X vssd1 vssd1 vccd1 vccd1 _13649_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15319_ _15333_/CLK _15319_/D vssd1 vssd1 vccd1 vccd1 _15319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16299_ _16312_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 _16299_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09811_ _15429_/Q _09867_/B _09811_/C vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__and3_1
XFILLER_99_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ _15419_/Q _09748_/C _09741_/X vssd1 vssd1 vccd1 vccd1 _09742_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09673_ _09671_/X _09672_/Y _09668_/B _09669_/C vssd1 vssd1 vccd1 vccd1 _09675_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _11229_/A vssd1 vssd1 vccd1 vccd1 _13051_/B sky130_fd_sc_hd__buf_6
XFILLER_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08555_ _15237_/Q _08560_/C _13045_/B vssd1 vssd1 vccd1 vccd1 _08557_/C sky130_fd_sc_hd__a21o_1
XFILLER_35_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08486_ _15228_/Q _08493_/C _13045_/B vssd1 vssd1 vccd1 vccd1 _08488_/C sky130_fd_sc_hd__a21o_1
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09107_ _09105_/Y _09100_/C _09102_/X _09103_/Y vssd1 vssd1 vccd1 vccd1 _09108_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09038_ _09038_/A vssd1 vssd1 vccd1 vccd1 _15308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11000_ _15615_/Q _11008_/C _10940_/X vssd1 vssd1 vccd1 vccd1 _11000_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12951_ _12949_/Y _12945_/C _12947_/X _12948_/Y vssd1 vssd1 vccd1 vccd1 _12952_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11902_ _12188_/A vssd1 vssd1 vccd1 vccd1 _11902_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15670_ _15763_/CLK _15670_/D vssd1 vssd1 vccd1 vccd1 _15670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12882_ _15911_/Q _12887_/C _12654_/X vssd1 vssd1 vccd1 vccd1 _12884_/C sky130_fd_sc_hd__a21o_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _16250_/Q _16249_/Q _16248_/Q _14620_/X vssd1 vssd1 vccd1 vccd1 _16233_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11833_ _15745_/Q _12007_/B _11833_/C vssd1 vssd1 vccd1 vccd1 _11843_/B sky130_fd_sc_hd__and3_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14552_/A _14552_/B _14552_/C vssd1 vssd1 vccd1 vccd1 _14553_/A sky130_fd_sc_hd__and3_1
X_11764_ _11762_/Y _11757_/C _11759_/X _11761_/Y vssd1 vssd1 vccd1 vccd1 _11765_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13604_/A _13503_/B _13507_/B vssd1 vssd1 vccd1 vccd1 _16013_/D sky130_fd_sc_hd__nor3_1
X_10715_ _15570_/Q _10722_/C _10655_/X vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _14482_/X _14481_/Y _14309_/X vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11695_ _15724_/Q _11811_/B _11697_/C vssd1 vssd1 vccd1 vccd1 _11695_/X sky130_fd_sc_hd__and3_1
X_16222_ _16222_/CLK _16222_/D vssd1 vssd1 vccd1 vccd1 _16222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ _13481_/A _13434_/B _13434_/C vssd1 vssd1 vccd1 vccd1 _13435_/A sky130_fd_sc_hd__and3_1
X_10646_ _11569_/A vssd1 vssd1 vccd1 vccd1 _10876_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16153_ _16166_/CLK _16153_/D vssd1 vssd1 vccd1 vccd1 _16153_/Q sky130_fd_sc_hd__dfxtp_2
X_13365_ _16007_/Q _16006_/Q _16005_/Q _13209_/X vssd1 vssd1 vccd1 vccd1 _15990_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_127_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10577_ _10577_/A _10577_/B _10577_/C vssd1 vssd1 vccd1 vccd1 _10579_/B sky130_fd_sc_hd__or3_1
XFILLER_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ _15110_/A _15103_/Y _15099_/B _15100_/C vssd1 vssd1 vccd1 vccd1 _15106_/B
+ sky130_fd_sc_hd__o211a_1
X_12316_ _12316_/A vssd1 vssd1 vccd1 vccd1 _15820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16084_ _16367_/CLK _16084_/D vssd1 vssd1 vccd1 vccd1 _16084_/Q sky130_fd_sc_hd__dfxtp_1
X_13296_ _13348_/A _13296_/B _13300_/B vssd1 vssd1 vccd1 vccd1 _15977_/D sky130_fd_sc_hd__nor3_1
XFILLER_142_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15035_ _15106_/A _15035_/B _15039_/B vssd1 vssd1 vccd1 vccd1 _16326_/D sky130_fd_sc_hd__nor3_1
X_12247_ _15817_/Q _15816_/Q _15815_/Q _12134_/X vssd1 vssd1 vccd1 vccd1 _15809_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12178_ _15799_/Q _12291_/B _12178_/C vssd1 vssd1 vccd1 vccd1 _12187_/B sky130_fd_sc_hd__and3_1
XFILLER_122_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11129_ _12277_/A vssd1 vssd1 vccd1 vccd1 _11362_/B sky130_fd_sc_hd__buf_2
XFILLER_96_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15937_ _15196_/Q _15937_/D vssd1 vssd1 vccd1 vccd1 _15937_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15868_ _15907_/CLK _15868_/D vssd1 vssd1 vccd1 vccd1 _15868_/Q sky130_fd_sc_hd__dfxtp_1
X_14819_ _16295_/Q _16294_/Q _16293_/Q _14818_/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__o31a_1
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15799_ _15195_/Q _15799_/D vssd1 vssd1 vccd1 vccd1 _15799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08340_ _08324_/A _08324_/B _08339_/X vssd1 vssd1 vccd1 vccd1 _08380_/B sky130_fd_sc_hd__o21ai_2
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08271_ _08271_/A _08271_/B vssd1 vssd1 vccd1 vccd1 _08272_/B sky130_fd_sc_hd__nor2_2
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07986_ _07986_/A _07888_/B vssd1 vssd1 vccd1 vccd1 _07986_/X sky130_fd_sc_hd__or2b_1
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09725_ _09746_/A _09725_/B _09725_/C vssd1 vssd1 vccd1 vccd1 _09726_/A sky130_fd_sc_hd__and3_1
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09656_ _15412_/Q _15411_/Q _15410_/Q _09541_/X vssd1 vssd1 vccd1 vccd1 _15404_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _08636_/C vssd1 vssd1 vccd1 vccd1 _08651_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09587_ _09594_/B _09587_/B vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__or2_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08538_ _08536_/A _08536_/B _08537_/X vssd1 vssd1 vccd1 vccd1 _15232_/D sky130_fd_sc_hd__a21oi_1
X_08469_ _08414_/X _08468_/Y _08466_/C _08421_/A vssd1 vssd1 vccd1 vccd1 _15222_/D
+ sky130_fd_sc_hd__a31oi_1
X_10500_ _15535_/Q _10729_/B _10506_/C vssd1 vssd1 vccd1 vccd1 _10500_/Y sky130_fd_sc_hd__nand3_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11480_ _15690_/Q _11487_/C _11425_/X vssd1 vssd1 vccd1 vccd1 _11480_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10431_ _10431_/A vssd1 vssd1 vccd1 vccd1 _15524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13150_ _13150_/A vssd1 vssd1 vccd1 vccd1 _15952_/D sky130_fd_sc_hd__clkbuf_1
X_10362_ _10362_/A vssd1 vssd1 vccd1 vccd1 _15514_/D sky130_fd_sc_hd__clkbuf_1
X_12101_ _15787_/Q _12102_/C _12100_/X vssd1 vssd1 vccd1 vccd1 _12101_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10293_ _15505_/Q _10331_/C _10181_/X vssd1 vssd1 vccd1 vccd1 _10297_/B sky130_fd_sc_hd__a21oi_1
X_13081_ _13081_/A _13081_/B vssd1 vssd1 vccd1 vccd1 _13082_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12032_ _12032_/A vssd1 vssd1 vccd1 vccd1 _15775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13983_ _16103_/Q _13990_/C _13982_/X vssd1 vssd1 vccd1 vccd1 _13985_/C sky130_fd_sc_hd__a21o_1
X_15722_ _15794_/CLK _15722_/D vssd1 vssd1 vccd1 vccd1 _15722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12934_ _12934_/A _12934_/B _12938_/A vssd1 vssd1 vccd1 vccd1 _15918_/D sky130_fd_sc_hd__nor3_1
X_15653_ _15655_/CLK _15653_/D vssd1 vssd1 vccd1 vccd1 _15653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12865_ _12865_/A _12865_/B vssd1 vssd1 vccd1 vccd1 _12869_/C sky130_fd_sc_hd__nor2_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14601_/B _14600_/Y _14601_/A vssd1 vssd1 vccd1 vccd1 _14604_/Y sky130_fd_sc_hd__o21bai_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _11814_/Y _11809_/C _11811_/X _11813_/Y vssd1 vssd1 vccd1 vccd1 _11817_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15584_/CLK _15584_/D vssd1 vssd1 vccd1 vccd1 _15584_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12796_/A _12796_/B _12796_/C vssd1 vssd1 vccd1 vccd1 _12797_/A sky130_fd_sc_hd__and3_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14368_/X _14533_/B _14528_/X vssd1 vssd1 vccd1 vccd1 _14535_/Y sky130_fd_sc_hd__a21oi_1
X_11747_ _11745_/X _11746_/Y _11742_/B _11743_/C vssd1 vssd1 vccd1 vccd1 _11749_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14466_ _16201_/Q _14546_/B _14466_/C vssd1 vssd1 vccd1 vccd1 _14471_/A sky130_fd_sc_hd__and3_1
X_11678_ _11697_/C vssd1 vssd1 vccd1 vccd1 _11712_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16205_ _16222_/CLK _16205_/D vssd1 vssd1 vccd1 vccd1 _16205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ _13430_/C vssd1 vssd1 vccd1 vccd1 _13445_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10629_ _10629_/A _10634_/C vssd1 vssd1 vccd1 vccd1 _10629_/X sky130_fd_sc_hd__or2_1
X_14397_ _14397_/A _14397_/B vssd1 vssd1 vccd1 vccd1 _14397_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16136_ _16148_/CLK _16136_/D vssd1 vssd1 vccd1 vccd1 _16136_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13348_ _13348_/A _13348_/B _13352_/B vssd1 vssd1 vccd1 vccd1 _15986_/D sky130_fd_sc_hd__nor3_1
XFILLER_6_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16067_ _16075_/CLK _16067_/D vssd1 vssd1 vccd1 vccd1 _16067_/Q sky130_fd_sc_hd__dfxtp_1
X_13279_ _13276_/X _13278_/Y _13272_/B _13273_/C vssd1 vssd1 vccd1 vccd1 _13281_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15018_ hold15/A _16339_/Q hold21/A _15017_/X vssd1 vssd1 vccd1 vccd1 _16323_/D sky130_fd_sc_hd__o31a_1
XFILLER_111_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07840_ _15917_/Q _15935_/Q vssd1 vssd1 vccd1 vccd1 _07842_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07771_ _15629_/Q _07771_/B _08069_/A vssd1 vssd1 vccd1 vccd1 _08069_/B sky130_fd_sc_hd__nand3_1
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09510_ _09508_/Y _09501_/C _09504_/X _09507_/Y vssd1 vssd1 vccd1 vccd1 _09511_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _09435_/B _09436_/C _09438_/X _09439_/Y vssd1 vssd1 vccd1 vccd1 _09442_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09372_ _15361_/Q _09372_/B _09380_/C vssd1 vssd1 vccd1 vccd1 _09377_/A sky130_fd_sc_hd__and3_1
XFILLER_40_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08323_ _08263_/A _08263_/B _08322_/Y vssd1 vssd1 vccd1 vccd1 _08324_/B sky130_fd_sc_hd__a21oi_2
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08254_ _08312_/A _08312_/B vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__xor2_4
XFILLER_118_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08185_ _07976_/A _07976_/B _08184_/X vssd1 vssd1 vccd1 vccd1 _08194_/A sky130_fd_sc_hd__o21ai_4
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07969_ _07969_/A vssd1 vssd1 vccd1 vccd1 _07973_/A sky130_fd_sc_hd__inv_2
X_09708_ _09708_/A _09708_/B _09708_/C vssd1 vssd1 vccd1 vccd1 _09710_/B sky130_fd_sc_hd__or3_1
XFILLER_56_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _10979_/B _10979_/C _10751_/X vssd1 vssd1 vccd1 vccd1 _10981_/C sky130_fd_sc_hd__o21ai_1
XFILLER_16_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _15402_/Q _09644_/C _09404_/X vssd1 vssd1 vccd1 vccd1 _09639_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12650_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12879_/B sky130_fd_sc_hd__buf_2
XFILLER_31_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11601_ _15707_/Q _11601_/B _11605_/C vssd1 vssd1 vccd1 vccd1 _11601_/Y sky130_fd_sc_hd__nand3_1
XFILLER_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12581_ _12579_/A _12579_/B _12580_/X vssd1 vssd1 vccd1 vccd1 _15861_/D sky130_fd_sc_hd__a21oi_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14320_ _14320_/A _14320_/B vssd1 vssd1 vccd1 vccd1 _14321_/B sky130_fd_sc_hd__and2_1
X_11532_ _11532_/A vssd1 vssd1 vccd1 vccd1 _15696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ _16157_/Q _14256_/C _14250_/X vssd1 vssd1 vccd1 vccd1 _14253_/C sky130_fd_sc_hd__a21o_1
XFILLER_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11463_ _15688_/Q _11525_/B _11466_/C vssd1 vssd1 vccd1 vccd1 _11463_/X sky130_fd_sc_hd__and3_1
XFILLER_99_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13202_ _13408_/A _13202_/B _13202_/C vssd1 vssd1 vccd1 vccd1 _13204_/B sky130_fd_sc_hd__or3_1
XFILLER_125_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10414_ _10446_/C vssd1 vssd1 vccd1 vccd1 _10453_/C sky130_fd_sc_hd__clkbuf_2
X_14182_ _14180_/A _14180_/B _14179_/Y _14181_/Y vssd1 vssd1 vccd1 vccd1 _16138_/D
+ sky130_fd_sc_hd__o31a_1
X_11394_ _11509_/A _11394_/B _11398_/A vssd1 vssd1 vccd1 vccd1 _15675_/D sky130_fd_sc_hd__nor3_1
XFILLER_125_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13133_ _15951_/Q _13293_/B _13138_/C vssd1 vssd1 vccd1 vccd1 _13133_/Y sky130_fd_sc_hd__nand3_1
XFILLER_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ _10345_/A vssd1 vssd1 vccd1 vccd1 _15511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _15942_/Q _13064_/B _13071_/C vssd1 vssd1 vccd1 vccd1 _13064_/X sky130_fd_sc_hd__and3_1
X_10276_ _15502_/Q _10512_/B _10276_/C vssd1 vssd1 vccd1 vccd1 _10284_/B sky130_fd_sc_hd__and3_1
XFILLER_140_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12015_ _12015_/A _12015_/B _12015_/C vssd1 vssd1 vccd1 vccd1 _12017_/B sky130_fd_sc_hd__or3_1
XFILLER_39_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13966_ _13921_/X _13964_/B _13922_/X vssd1 vssd1 vccd1 vccd1 _13966_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15705_ _15794_/CLK _15705_/D vssd1 vssd1 vccd1 vccd1 _15705_/Q sky130_fd_sc_hd__dfxtp_1
X_12917_ _12917_/A _12917_/B vssd1 vssd1 vccd1 vccd1 _12918_/B sky130_fd_sc_hd__nor2_1
X_13897_ _14414_/A vssd1 vssd1 vccd1 vccd1 _14883_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15636_ _15194_/Q _15636_/D vssd1 vssd1 vccd1 vccd1 _15636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12848_ _15904_/Q _13066_/B _12854_/C vssd1 vssd1 vccd1 vccd1 _12848_/Y sky130_fd_sc_hd__nand3_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15567_ _15655_/CLK _15567_/D vssd1 vssd1 vccd1 vccd1 _15567_/Q sky130_fd_sc_hd__dfxtp_2
X_12779_ _15894_/Q _12786_/C _12661_/X vssd1 vssd1 vccd1 vccd1 _12779_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _16213_/Q _14598_/B _14525_/C vssd1 vssd1 vccd1 vccd1 _14521_/A sky130_fd_sc_hd__and3_1
X_15498_ _15224_/Q _15498_/D vssd1 vssd1 vccd1 vccd1 _15498_/Q sky130_fd_sc_hd__dfxtp_1
X_14449_ _14447_/X _14449_/B vssd1 vssd1 vccd1 vccd1 _14449_/X sky130_fd_sc_hd__and2b_1
XFILLER_116_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16119_ _16119_/CLK _16119_/D vssd1 vssd1 vccd1 vccd1 _16119_/Q sky130_fd_sc_hd__dfxtp_1
X_09990_ _15457_/Q _09989_/C _09755_/X vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__a21oi_1
X_08941_ _08939_/Y _08934_/C _08937_/X _08938_/Y vssd1 vssd1 vccd1 vccd1 _08942_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_97_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08872_ _15285_/Q _08872_/B _08880_/C vssd1 vssd1 vccd1 vccd1 _08872_/X sky130_fd_sc_hd__and3_1
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07823_ _08044_/A _07823_/B vssd1 vssd1 vccd1 vccd1 _07825_/B sky130_fd_sc_hd__xnor2_2
XFILLER_69_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07754_ _15954_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07755_/B sky130_fd_sc_hd__or2_1
XFILLER_53_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07685_ _14806_/A vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_91_clk _15584_/CLK vssd1 vssd1 vccd1 vccd1 _15602_/CLK sky130_fd_sc_hd__clkbuf_16
X_09424_ _15368_/Q vssd1 vssd1 vccd1 vccd1 _09438_/C sky130_fd_sc_hd__inv_2
XFILLER_52_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09355_ _15359_/Q _09354_/C _09180_/X vssd1 vssd1 vccd1 vccd1 _09356_/B sky130_fd_sc_hd__a21oi_1
XFILLER_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ _08306_/A _08239_/A vssd1 vssd1 vccd1 vccd1 _08306_/X sky130_fd_sc_hd__or2b_1
X_09286_ _09283_/X _09284_/Y _09285_/Y _09281_/C vssd1 vssd1 vccd1 vccd1 _09288_/B
+ sky130_fd_sc_hd__o211ai_1
X_08237_ _08115_/A _08115_/B _08236_/X vssd1 vssd1 vccd1 vccd1 _08238_/B sky130_fd_sc_hd__a21oi_2
XFILLER_4_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08168_ _14316_/A vssd1 vssd1 vccd1 vccd1 _08168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08099_ _08099_/A vssd1 vssd1 vccd1 vccd1 _14863_/C sky130_fd_sc_hd__clkbuf_2
X_10130_ _10131_/B _10131_/C _10131_/A vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__a21o_1
XFILLER_121_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10061_ _10100_/C vssd1 vssd1 vccd1 vccd1 _10106_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13820_ _13832_/C vssd1 vssd1 vccd1 vccd1 _13846_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ _13868_/A vssd1 vssd1 vccd1 vccd1 _13852_/A sky130_fd_sc_hd__buf_2
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10963_ _15609_/Q _10963_/B _10963_/C vssd1 vssd1 vccd1 vccd1 _10973_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_82_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15440_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12702_ _12702_/A vssd1 vssd1 vccd1 vccd1 _15880_/D sky130_fd_sc_hd__clkbuf_1
X_13682_ _13683_/B _13683_/C _13683_/A vssd1 vssd1 vccd1 vccd1 _13684_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10894_ _10894_/A vssd1 vssd1 vccd1 vccd1 _15597_/D sky130_fd_sc_hd__clkbuf_1
X_15421_ _15484_/CLK _15421_/D vssd1 vssd1 vccd1 vccd1 _15421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12633_ _12640_/B _12633_/B vssd1 vssd1 vccd1 vccd1 _12635_/A sky130_fd_sc_hd__or2_1
XFILLER_43_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16376__25 vssd1 vssd1 vccd1 vccd1 _16376__25/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15352_ _15368_/CLK _15352_/D vssd1 vssd1 vccd1 vccd1 _15352_/Q sky130_fd_sc_hd__dfxtp_2
X_12564_ _12562_/Y _12557_/C _12559_/X _12560_/Y vssd1 vssd1 vccd1 vccd1 _12565_/C
+ sky130_fd_sc_hd__a211o_1
X_14303_ _14295_/B _14296_/C _14307_/A _14301_/Y vssd1 vssd1 vccd1 vccd1 _14307_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11515_ _11515_/A _11515_/B _11515_/C vssd1 vssd1 vccd1 vccd1 _11516_/C sky130_fd_sc_hd__nand3_1
XFILLER_12_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15283_ _15301_/CLK _15283_/D vssd1 vssd1 vccd1 vccd1 _15283_/Q sky130_fd_sc_hd__dfxtp_1
X_12495_ _12488_/B _12489_/C _12492_/X _12493_/Y vssd1 vssd1 vccd1 vccd1 _12496_/C
+ sky130_fd_sc_hd__a211o_1
X_14234_ _14320_/A _14234_/B vssd1 vssd1 vccd1 vccd1 _14235_/B sky130_fd_sc_hd__and2_1
X_11446_ _11466_/C vssd1 vssd1 vccd1 vccd1 _11479_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14165_ _16139_/Q _14249_/B _14171_/C vssd1 vssd1 vccd1 vccd1 _14168_/B sky130_fd_sc_hd__nand3_1
X_11377_ _11377_/A _11377_/B vssd1 vssd1 vccd1 vccd1 _11378_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ _13640_/A vssd1 vssd1 vccd1 vccd1 _13333_/B sky130_fd_sc_hd__buf_2
X_10328_ _10336_/A _10326_/Y _10327_/Y _10323_/C vssd1 vssd1 vccd1 vccd1 _10330_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _14102_/A _14094_/Y _14095_/Y _14091_/C vssd1 vssd1 vccd1 vccd1 _14098_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13048_/B _13048_/C _13048_/A vssd1 vssd1 vccd1 vccd1 _13049_/B sky130_fd_sc_hd__a21o_1
X_10259_ _10266_/A _10259_/B _10259_/C vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__and3_1
XFILLER_140_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14998_ _14998_/A _14998_/B vssd1 vssd1 vccd1 vccd1 _14999_/B sky130_fd_sc_hd__nor2_1
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13949_ _13980_/A _13949_/B _13952_/B vssd1 vssd1 vccd1 vccd1 _16092_/D sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_73_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15333_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ _15194_/Q _15619_/D vssd1 vssd1 vccd1 vccd1 _15619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09140_ _09160_/C vssd1 vssd1 vccd1 vccd1 _09173_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09071_ _09071_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09075_/C sky130_fd_sc_hd__nor2_1
X_08022_ _15854_/Q _08022_/B vssd1 vssd1 vccd1 vccd1 _08022_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09973_ _15455_/Q _09979_/C _09741_/X vssd1 vssd1 vccd1 vccd1 _09973_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08924_ _08942_/A _08924_/B _08924_/C vssd1 vssd1 vccd1 vccd1 _08925_/A sky130_fd_sc_hd__and3_1
XFILLER_130_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08855_ _08856_/B _08856_/C _08856_/A vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__a21o_1
XFILLER_111_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07806_ _14289_/C _07807_/B vssd1 vssd1 vccd1 vccd1 _07808_/A sky130_fd_sc_hd__nand2_1
XFILLER_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08786_ _08786_/A vssd1 vssd1 vccd1 vccd1 _15269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07737_ _07737_/A vssd1 vssd1 vccd1 vccd1 _15024_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_64_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16353_/CLK sky130_fd_sc_hd__clkbuf_16
X_07668_ _15030_/A _07668_/B vssd1 vssd1 vccd1 vccd1 _07668_/X sky130_fd_sc_hd__or2_1
XFILLER_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09407_ _09414_/A _09405_/Y _09406_/Y _09401_/C vssd1 vssd1 vccd1 vccd1 _09409_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07599_ _14459_/A vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09338_ _09338_/A vssd1 vssd1 vccd1 vccd1 _15355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ _10134_/A vssd1 vssd1 vccd1 vccd1 _09496_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11300_ _11298_/Y _11293_/C _11296_/X _11297_/Y vssd1 vssd1 vccd1 vccd1 _11301_/C
+ sky130_fd_sc_hd__a211o_1
X_12280_ _12278_/Y _12273_/C _12275_/X _12276_/Y vssd1 vssd1 vccd1 vccd1 _12281_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11231_ _15651_/Q _11239_/C _11230_/X vssd1 vssd1 vccd1 vccd1 _11231_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11162_ _11220_/A _11162_/B _11166_/A vssd1 vssd1 vccd1 vccd1 _15639_/D sky130_fd_sc_hd__nor3_1
XFILLER_107_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10113_ _10111_/A _10111_/B _10112_/X vssd1 vssd1 vccd1 vccd1 _15474_/D sky130_fd_sc_hd__a21oi_1
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11093_ _11267_/A vssd1 vssd1 vccd1 vccd1 _11133_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15970_ _15970_/CLK _15970_/D vssd1 vssd1 vccd1 vccd1 _15970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10044_ _10044_/A vssd1 vssd1 vccd1 vccd1 _10044_/X sky130_fd_sc_hd__clkbuf_2
X_14921_ _14921_/A _14921_/B vssd1 vssd1 vccd1 vccd1 _14922_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14852_ _15050_/A vssd1 vssd1 vccd1 vccd1 _15010_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13803_ _13801_/Y _13797_/C _13808_/A _13800_/Y vssd1 vssd1 vccd1 vccd1 _13808_/B
+ sky130_fd_sc_hd__a211oi_1
X_14783_ hold12/A _14782_/C _14744_/X vssd1 vssd1 vccd1 vccd1 _14785_/C sky130_fd_sc_hd__a21o_1
X_11995_ _11991_/X _11992_/Y _11994_/Y _11989_/C vssd1 vssd1 vccd1 vccd1 _11997_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_91_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _16312_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13734_ _13734_/A _13734_/B _13734_/C vssd1 vssd1 vccd1 vccd1 _13735_/C sky130_fd_sc_hd__nand3_1
X_10946_ _15607_/Q _10950_/B _11128_/A vssd1 vssd1 vccd1 vccd1 _10946_/X sky130_fd_sc_hd__and3_1
XFILLER_71_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13665_ _13665_/A vssd1 vssd1 vccd1 vccd1 _16042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10877_ _15596_/Q _10882_/C _10648_/X vssd1 vssd1 vccd1 vccd1 _10879_/C sky130_fd_sc_hd__a21o_1
X_15404_ _15422_/CLK _15404_/D vssd1 vssd1 vccd1 vccd1 _15404_/Q sky130_fd_sc_hd__dfxtp_1
X_12616_ _12616_/A vssd1 vssd1 vccd1 vccd1 _12616_/X sky130_fd_sc_hd__buf_2
X_13596_ _13596_/A vssd1 vssd1 vccd1 vccd1 _16030_/D sky130_fd_sc_hd__clkbuf_1
X_15335_ _15337_/CLK _15335_/D vssd1 vssd1 vccd1 vccd1 _15335_/Q sky130_fd_sc_hd__dfxtp_1
X_12547_ _15858_/Q _12554_/C _12377_/X vssd1 vssd1 vccd1 vccd1 _12547_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_145_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15266_ _15274_/CLK _15266_/D vssd1 vssd1 vccd1 vccd1 _15266_/Q sky130_fd_sc_hd__dfxtp_1
X_12478_ _12492_/C vssd1 vssd1 vccd1 vccd1 _12500_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_3 state1[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ _16149_/Q _14216_/C _14033_/X vssd1 vssd1 vccd1 vccd1 _14217_/Y sky130_fd_sc_hd__a21oi_1
X_11429_ _11427_/Y _11420_/C _11434_/A _11426_/Y vssd1 vssd1 vccd1 vccd1 _11434_/B
+ sky130_fd_sc_hd__a211oi_1
X_15197_ _16353_/CLK _15197_/D vssd1 vssd1 vccd1 vccd1 spike_out[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_99_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14148_ _14328_/A vssd1 vssd1 vccd1 vccd1 _14368_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14079_ _14079_/A vssd1 vssd1 vccd1 vccd1 _16118_/D sky130_fd_sc_hd__clkbuf_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08640_ _08640_/A vssd1 vssd1 vccd1 vccd1 _15247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ _08580_/A _08571_/B _08571_/C vssd1 vssd1 vccd1 vccd1 _08572_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_46_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _16247_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09123_ _09202_/A _09123_/B _09128_/B vssd1 vssd1 vccd1 vccd1 _15321_/D sky130_fd_sc_hd__nor3_1
XFILLER_148_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09054_ _13693_/A vssd1 vssd1 vccd1 vccd1 _09285_/B sky130_fd_sc_hd__buf_2
X_08005_ _15963_/Q vssd1 vssd1 vccd1 vccd1 _13266_/C sky130_fd_sc_hd__inv_2
XFILLER_144_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _09977_/A _09956_/B _09956_/C vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__and3_1
XFILLER_106_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08907_ _15290_/Q _08951_/C _08735_/X vssd1 vssd1 vccd1 vccd1 _08909_/B sky130_fd_sc_hd__a21oi_1
X_09887_ _09887_/A vssd1 vssd1 vccd1 vccd1 _15439_/D sky130_fd_sc_hd__clkbuf_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08838_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08878_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08769_ _15268_/Q _09001_/B _08769_/C vssd1 vssd1 vccd1 vccd1 _08778_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_37_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _16222_/CLK sky130_fd_sc_hd__clkbuf_16
X_10800_ _10806_/B _10800_/B vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__or2_1
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11780_ _11780_/A _11784_/C vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__or2_1
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10731_ _10729_/Y _10725_/C _10727_/X _10728_/Y vssd1 vssd1 vccd1 vccd1 _10732_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13450_ _13476_/A _13450_/B _13455_/B vssd1 vssd1 vccd1 vccd1 _16004_/D sky130_fd_sc_hd__nor3_1
X_10662_ _15562_/Q _10888_/B _10665_/C vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__and3_1
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12401_ _15833_/Q _12458_/B _12405_/C vssd1 vssd1 vccd1 vccd1 _12401_/Y sky130_fd_sc_hd__nand3_1
XFILLER_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13381_ _15995_/Q _13380_/C _13277_/X vssd1 vssd1 vccd1 vccd1 _13381_/Y sky130_fd_sc_hd__a21oi_1
X_10593_ _10593_/A _10593_/B _10593_/C vssd1 vssd1 vccd1 vccd1 _10594_/C sky130_fd_sc_hd__nand3_1
X_15120_ _15189_/A _15189_/B _15120_/C vssd1 vssd1 vccd1 vccd1 _15122_/A sky130_fd_sc_hd__and3_1
X_12332_ _12616_/A vssd1 vssd1 vccd1 vccd1 _12332_/X sky130_fd_sc_hd__buf_2
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15051_ _15051_/A _15189_/B _15051_/C vssd1 vssd1 vccd1 vccd1 _15053_/A sky130_fd_sc_hd__and3_1
X_12263_ _15813_/Q _12270_/C _12093_/X vssd1 vssd1 vccd1 vccd1 _12263_/Y sky130_fd_sc_hd__a21oi_1
X_14002_ _13999_/B _13998_/Y _13999_/A vssd1 vssd1 vccd1 vccd1 _14002_/Y sky130_fd_sc_hd__o21bai_1
X_11214_ _11228_/C vssd1 vssd1 vccd1 vccd1 _11239_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12194_ _12208_/C vssd1 vssd1 vccd1 vccd1 _12216_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11145_ _11151_/B _11145_/B vssd1 vssd1 vccd1 vccd1 _11147_/A sky130_fd_sc_hd__or2_1
XFILLER_96_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11076_ _11076_/A _11076_/B _11076_/C vssd1 vssd1 vccd1 vccd1 _11077_/A sky130_fd_sc_hd__and3_1
X_15953_ _15970_/CLK _15953_/D vssd1 vssd1 vccd1 vccd1 _15953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10027_ _10035_/A _10027_/B _10027_/C vssd1 vssd1 vccd1 vccd1 _10028_/A sky130_fd_sc_hd__and3_1
X_14904_ _14915_/A _14904_/B _14908_/A vssd1 vssd1 vccd1 vccd1 _16297_/D sky130_fd_sc_hd__nor3_1
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15884_ _07603_/A _15884_/D vssd1 vssd1 vccd1 vccd1 _15884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14835_ _14841_/A _14834_/Y _14829_/B _14830_/C vssd1 vssd1 vccd1 vccd1 _14837_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_clk clkbuf_3_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15970_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11978_ _15768_/Q _12150_/B _11978_/C vssd1 vssd1 vccd1 vccd1 _11978_/X sky130_fd_sc_hd__and3_1
X_14766_ _14964_/A vssd1 vssd1 vccd1 vccd1 _14766_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10929_ _15604_/Q _10970_/B _10760_/X vssd1 vssd1 vccd1 vccd1 _10931_/B sky130_fd_sc_hd__a21oi_1
X_13717_ _13716_/B _13716_/C _13562_/X vssd1 vssd1 vccd1 vccd1 _13718_/C sky130_fd_sc_hd__o21ai_1
X_14697_ _14697_/A _14697_/B vssd1 vssd1 vccd1 vccd1 _16249_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13648_ _16042_/Q _13648_/B _13648_/C vssd1 vssd1 vccd1 vccd1 _13658_/A sky130_fd_sc_hd__and3_1
XFILLER_20_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13579_ _13580_/B _13580_/C _13580_/A vssd1 vssd1 vccd1 vccd1 _13581_/B sky130_fd_sc_hd__a21o_1
X_16367_ _16367_/CLK _16367_/D vssd1 vssd1 vccd1 vccd1 _16367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15318_ _15333_/CLK _15318_/D vssd1 vssd1 vccd1 vccd1 _15318_/Q sky130_fd_sc_hd__dfxtp_1
X_16298_ _16312_/CLK _16298_/D vssd1 vssd1 vccd1 vccd1 _16298_/Q sky130_fd_sc_hd__dfxtp_2
X_15249_ _15259_/CLK _15249_/D vssd1 vssd1 vccd1 vccd1 _15249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09810_ _10388_/A vssd1 vssd1 vccd1 vccd1 _09930_/A sky130_fd_sc_hd__buf_2
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09741_ _10610_/A vssd1 vssd1 vccd1 vccd1 _09741_/X sky130_fd_sc_hd__clkbuf_2
X_09672_ _15408_/Q _09680_/C _09497_/X vssd1 vssd1 vccd1 vccd1 _09672_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08623_ input3/X vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__buf_2
XFILLER_94_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _15984_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _15237_/Q _13526_/A _08560_/C vssd1 vssd1 vccd1 vccd1 _08557_/B sky130_fd_sc_hd__nand3_1
XFILLER_70_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08485_ _15228_/Q _13526_/A _08493_/C vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__nand3_1
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09106_ _09102_/X _09103_/Y _09105_/Y _09100_/C vssd1 vssd1 vccd1 vccd1 _09108_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_109_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09037_ _09058_/A _09037_/B _09037_/C vssd1 vssd1 vccd1 vccd1 _09038_/A sky130_fd_sc_hd__and3_1
XFILLER_108_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09939_ _09997_/A _09939_/B _09939_/C vssd1 vssd1 vccd1 vccd1 _09941_/B sky130_fd_sc_hd__or3_1
X_12950_ _12947_/X _12948_/Y _12949_/Y _12945_/C vssd1 vssd1 vccd1 vccd1 _12952_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11901_ _12015_/A _11901_/B _11901_/C vssd1 vssd1 vccd1 vccd1 _11904_/B sky130_fd_sc_hd__or3_1
X_12881_ _15911_/Q _12935_/B _12887_/C vssd1 vssd1 vccd1 vccd1 _12884_/B sky130_fd_sc_hd__nand3_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11832_ _11949_/A _11832_/B _11836_/B vssd1 vssd1 vccd1 vccd1 _15743_/D sky130_fd_sc_hd__nor3_1
X_14620_ _14818_/A vssd1 vssd1 vccd1 vccd1 _14620_/X sky130_fd_sc_hd__buf_2
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14551_/A _14551_/B _14551_/C vssd1 vssd1 vccd1 vccd1 _14552_/C sky130_fd_sc_hd__nand3_1
X_11763_ _11759_/X _11761_/Y _11762_/Y _11757_/C vssd1 vssd1 vccd1 vccd1 _11765_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _15570_/Q _10999_/B _10714_/C vssd1 vssd1 vccd1 vccd1 _10714_/X sky130_fd_sc_hd__and3_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13500_/Y _13495_/C _13507_/A _13499_/Y vssd1 vssd1 vccd1 vccd1 _13507_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14482_/A _14482_/B vssd1 vssd1 vccd1 vccd1 _14482_/X sky130_fd_sc_hd__or2_1
X_11694_ _11694_/A vssd1 vssd1 vccd1 vccd1 _15722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16221_ _16362_/CLK _16221_/D vssd1 vssd1 vccd1 vccd1 _16221_/Q sky130_fd_sc_hd__dfxtp_1
X_13433_ _13427_/B _13428_/C _13430_/X _13431_/Y vssd1 vssd1 vccd1 vccd1 _13434_/C
+ sky130_fd_sc_hd__a211o_1
X_10645_ _10645_/A _10645_/B _10651_/A vssd1 vssd1 vccd1 vccd1 _15558_/D sky130_fd_sc_hd__nor3_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16152_ _16187_/CLK _16152_/D vssd1 vssd1 vccd1 vccd1 _16152_/Q sky130_fd_sc_hd__dfxtp_1
X_13364_ _13153_/X _13360_/C _13363_/Y vssd1 vssd1 vccd1 vccd1 _15989_/D sky130_fd_sc_hd__a21oi_1
X_10576_ _10693_/A vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15103_ _16348_/Q _15107_/C _14988_/X vssd1 vssd1 vccd1 vccd1 _15103_/Y sky130_fd_sc_hd__a21oi_1
X_12315_ _12337_/A _12315_/B _12315_/C vssd1 vssd1 vccd1 vccd1 _12316_/A sky130_fd_sc_hd__and3_1
X_16083_ _16367_/CLK _16083_/D vssd1 vssd1 vccd1 vccd1 _16083_/Q sky130_fd_sc_hd__dfxtp_2
X_13295_ _13293_/Y _13289_/C _13300_/A _13292_/Y vssd1 vssd1 vccd1 vccd1 _13300_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _15027_/B _15028_/C _15039_/A _15032_/Y vssd1 vssd1 vccd1 vccd1 _15039_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12246_ _12246_/A vssd1 vssd1 vccd1 vccd1 _15808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12177_ _12234_/A _12177_/B _12181_/B vssd1 vssd1 vccd1 vccd1 _15797_/D sky130_fd_sc_hd__nor3_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _11128_/A vssd1 vssd1 vccd1 vccd1 _12277_/A sky130_fd_sc_hd__buf_4
XFILLER_68_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11059_ _15624_/Q _11066_/C _10940_/X vssd1 vssd1 vccd1 vccd1 _11059_/Y sky130_fd_sc_hd__a21oi_1
X_15936_ _16100_/CLK _15936_/D vssd1 vssd1 vccd1 vccd1 _15936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15867_ _07603_/A _15867_/D vssd1 vssd1 vccd1 vccd1 _15867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14818_ _14818_/A vssd1 vssd1 vccd1 vccd1 _14818_/X sky130_fd_sc_hd__buf_2
X_15798_ _15195_/Q _15798_/D vssd1 vssd1 vccd1 vccd1 _15798_/Q sky130_fd_sc_hd__dfxtp_1
X_14749_ _14749_/A vssd1 vssd1 vccd1 vccd1 _16262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08270_ _08270_/A _08270_/B _08270_/C vssd1 vssd1 vccd1 vccd1 _08271_/B sky130_fd_sc_hd__and3_1
XFILLER_149_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_opt_3_0_clk clkbuf_3_4_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clk _15818_/CLK vssd1 vssd1 vccd1 vccd1 _15809_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07985_ _08178_/A _07985_/B vssd1 vssd1 vccd1 vccd1 _08151_/A sky130_fd_sc_hd__xnor2_4
X_09724_ _09724_/A _09724_/B _09724_/C vssd1 vssd1 vccd1 vccd1 _09725_/C sky130_fd_sc_hd__nand3_1
XFILLER_68_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ _09655_/A vssd1 vssd1 vccd1 vccd1 _15403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08606_ _08622_/C vssd1 vssd1 vccd1 vccd1 _08636_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09586_ _15394_/Q _09585_/C _09467_/X vssd1 vssd1 vccd1 vccd1 _09587_/B sky130_fd_sc_hd__a21oi_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 _15818_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _15030_/A _08540_/C vssd1 vssd1 vccd1 vccd1 _08537_/X sky130_fd_sc_hd__or2_1
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08468_ _08468_/A _08468_/B vssd1 vssd1 vccd1 vccd1 _08468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08399_ _08411_/A _08397_/Y _08372_/A _08378_/A vssd1 vssd1 vccd1 vccd1 _08400_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_10_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ _10444_/A _10430_/B _10430_/C vssd1 vssd1 vccd1 vccd1 _10431_/A sky130_fd_sc_hd__and3_1
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10361_ _10386_/A _10361_/B _10361_/C vssd1 vssd1 vccd1 vccd1 _10362_/A sky130_fd_sc_hd__and3_1
X_12100_ _12100_/A vssd1 vssd1 vccd1 vccd1 _12100_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13080_ _13086_/B _13080_/B vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__or2_1
X_10292_ _10325_/C vssd1 vssd1 vccd1 vccd1 _10331_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_88_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _12053_/A _12031_/B _12031_/C vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__and3_1
XFILLER_88_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13982_ _14250_/A vssd1 vssd1 vccd1 vccd1 _13982_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15721_ _15794_/CLK _15721_/D vssd1 vssd1 vccd1 vccd1 _15721_/Q sky130_fd_sc_hd__dfxtp_1
X_12933_ _15919_/Q _13043_/B _12941_/C vssd1 vssd1 vccd1 vccd1 _12938_/A sky130_fd_sc_hd__and3_1
XFILLER_37_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15652_ _15655_/CLK _15652_/D vssd1 vssd1 vccd1 vccd1 _15652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12864_/A _12864_/B vssd1 vssd1 vccd1 vccd1 _12865_/B sky130_fd_sc_hd__nor2_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14601_/A _14601_/B _14600_/Y _14602_/Y vssd1 vssd1 vccd1 vccd1 _16228_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _11811_/X _11813_/Y _11814_/Y _11809_/C vssd1 vssd1 vccd1 vccd1 _11817_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _15655_/CLK _15583_/D vssd1 vssd1 vccd1 vccd1 _15583_/Q sky130_fd_sc_hd__dfxtp_1
X_12795_ _12793_/Y _12789_/C _12791_/X _12792_/Y vssd1 vssd1 vccd1 vccd1 _12796_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _15732_/Q _11754_/C _11519_/X vssd1 vssd1 vccd1 vccd1 _11746_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14534_ _14408_/X _14532_/B _14533_/Y vssd1 vssd1 vccd1 vccd1 _16212_/D sky130_fd_sc_hd__o21a_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11677_ _11689_/C vssd1 vssd1 vccd1 vccd1 _11697_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14465_ _16201_/Q _14486_/C _14287_/X vssd1 vssd1 vccd1 vccd1 _14467_/B sky130_fd_sc_hd__a21oi_1
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16204_ _16204_/CLK _16204_/D vssd1 vssd1 vccd1 vccd1 _16204_/Q sky130_fd_sc_hd__dfxtp_1
X_10628_ _10628_/A _10628_/B vssd1 vssd1 vccd1 vccd1 _10634_/C sky130_fd_sc_hd__nor2_1
X_13416_ _13420_/C vssd1 vssd1 vccd1 vccd1 _13430_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14396_ _16186_/Q _14403_/C _14395_/X vssd1 vssd1 vccd1 vccd1 _14398_/B sky130_fd_sc_hd__a21oi_1
XFILLER_127_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13347_ _13345_/Y _13339_/C _13352_/A _13343_/Y vssd1 vssd1 vccd1 vccd1 _13352_/B
+ sky130_fd_sc_hd__a211oi_1
X_16135_ _16148_/CLK _16135_/D vssd1 vssd1 vccd1 vccd1 _16135_/Q sky130_fd_sc_hd__dfxtp_2
X_10559_ _10559_/A _10559_/B _10559_/C vssd1 vssd1 vccd1 vccd1 _10560_/A sky130_fd_sc_hd__and3_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16066_ _16075_/CLK _16066_/D vssd1 vssd1 vccd1 vccd1 _16066_/Q sky130_fd_sc_hd__dfxtp_1
X_13278_ _15977_/Q _13276_/C _13277_/X vssd1 vssd1 vccd1 vccd1 _13278_/Y sky130_fd_sc_hd__a21oi_1
X_12229_ _15807_/Q _12235_/C _12001_/X vssd1 vssd1 vccd1 vccd1 _12229_/Y sky130_fd_sc_hd__a21oi_1
X_15017_ _15017_/A vssd1 vssd1 vccd1 vccd1 _15017_/X sky130_fd_sc_hd__buf_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07770_ _07771_/B _08069_/A _15629_/Q vssd1 vssd1 vccd1 vccd1 _07772_/A sky130_fd_sc_hd__a21o_1
XFILLER_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15919_ _15196_/Q _15919_/D vssd1 vssd1 vccd1 vccd1 _15919_/Q sky130_fd_sc_hd__dfxtp_1
X_09440_ _09438_/X _09439_/Y _09435_/B _09436_/C vssd1 vssd1 vccd1 vccd1 _09442_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09371_ _15361_/Q _09411_/C _09316_/X vssd1 vssd1 vccd1 vccd1 _09373_/B sky130_fd_sc_hd__a21oi_1
XFILLER_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08322_ _08322_/A _08322_/B vssd1 vssd1 vccd1 vccd1 _08322_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08253_ _08139_/A _08139_/B _08252_/Y vssd1 vssd1 vccd1 vccd1 _08312_/B sky130_fd_sc_hd__a21oi_2
X_08184_ _08184_/A _07977_/A vssd1 vssd1 vccd1 vccd1 _08184_/X sky130_fd_sc_hd__or2b_1
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07968_ _14426_/C _14505_/C _07967_/Y vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__o21ai_1
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09707_ _09825_/A vssd1 vssd1 vccd1 vccd1 _09746_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07899_ _15584_/Q vssd1 vssd1 vccd1 vccd1 _10812_/A sky130_fd_sc_hd__clkinv_2
XFILLER_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09638_ _15402_/Q _09867_/B _09638_/C vssd1 vssd1 vccd1 vccd1 _09647_/A sky130_fd_sc_hd__and3_1
XFILLER_71_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09569_ _09569_/A vssd1 vssd1 vccd1 vccd1 _15390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11600_ _15708_/Q _11605_/C _11425_/X vssd1 vssd1 vccd1 vccd1 _11600_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _12636_/A _12583_/C vssd1 vssd1 vccd1 vccd1 _12580_/X sky130_fd_sc_hd__or2_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11531_ _11538_/A _11531_/B _11531_/C vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__and3_1
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _14250_/A vssd1 vssd1 vccd1 vccd1 _14250_/X sky130_fd_sc_hd__clkbuf_4
X_11462_ _11462_/A vssd1 vssd1 vccd1 vccd1 _15686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _15050_/A vssd1 vssd1 vccd1 vccd1 _13408_/A sky130_fd_sc_hd__clkbuf_2
X_10413_ _10434_/C vssd1 vssd1 vccd1 vccd1 _10446_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14181_ _14180_/X _14179_/Y _14042_/X vssd1 vssd1 vccd1 vccd1 _14181_/Y sky130_fd_sc_hd__a21oi_1
X_11393_ _15676_/Q _11449_/B _11401_/C vssd1 vssd1 vccd1 vccd1 _11398_/A sky130_fd_sc_hd__and3_1
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ _14395_/A vssd1 vssd1 vccd1 vccd1 _13293_/B sky130_fd_sc_hd__buf_4
X_10344_ _10386_/A _10344_/B _10344_/C vssd1 vssd1 vccd1 vccd1 _10345_/A sky130_fd_sc_hd__and3_1
XFILLER_124_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13063_ _13063_/A vssd1 vssd1 vccd1 vccd1 _15940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10275_ _11197_/A vssd1 vssd1 vccd1 vccd1 _10512_/B sky130_fd_sc_hd__clkbuf_2
X_12014_ _12129_/A vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13965_ _13912_/X _13963_/B _13964_/Y vssd1 vssd1 vccd1 vccd1 _16095_/D sky130_fd_sc_hd__o21a_1
X_15704_ _15794_/CLK _15704_/D vssd1 vssd1 vccd1 vccd1 _15704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12916_ _12923_/B _12916_/B vssd1 vssd1 vccd1 vccd1 _12918_/A sky130_fd_sc_hd__or2_1
X_13896_ _13896_/A _13896_/B vssd1 vssd1 vccd1 vccd1 _13896_/X sky130_fd_sc_hd__or2_1
XFILLER_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15635_ _15194_/Q _15635_/D vssd1 vssd1 vccd1 vccd1 _15635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12847_/A vssd1 vssd1 vccd1 vccd1 _13066_/B sky130_fd_sc_hd__buf_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15566_ _15575_/CLK _15566_/D vssd1 vssd1 vccd1 vccd1 _15566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _15894_/Q _12996_/B _12778_/C vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__and3_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14517_ _14517_/A _14517_/B _14520_/B vssd1 vssd1 vccd1 vccd1 _16209_/D sky130_fd_sc_hd__nor3_1
X_11729_ _11765_/A _11729_/B _11729_/C vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__and3_1
XFILLER_30_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15497_ _15224_/Q _15497_/D vssd1 vssd1 vccd1 vccd1 _15497_/Q sky130_fd_sc_hd__dfxtp_1
X_14448_ _16196_/Q _14447_/C _14270_/X vssd1 vssd1 vccd1 vccd1 _14449_/B sky130_fd_sc_hd__a21o_1
XFILLER_116_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14379_ _14379_/A vssd1 vssd1 vccd1 vccd1 _14546_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_128_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16118_ _16129_/CLK _16118_/D vssd1 vssd1 vccd1 vccd1 _16118_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16049_ _16050_/CLK _16049_/D vssd1 vssd1 vccd1 vccd1 _16049_/Q sky130_fd_sc_hd__dfxtp_1
X_08940_ _08937_/X _08938_/Y _08939_/Y _08934_/C vssd1 vssd1 vccd1 vccd1 _08942_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_103_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08871_ _08871_/A vssd1 vssd1 vccd1 vccd1 _15283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07822_ _07822_/A _07822_/B vssd1 vssd1 vccd1 vccd1 _07823_/B sky130_fd_sc_hd__xor2_2
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07753_ _15954_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07755_/A sky130_fd_sc_hd__nand2_1
X_07684_ _14364_/A vssd1 vssd1 vccd1 vccd1 _14806_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ _15376_/Q _15375_/Q _15374_/Q _09194_/X vssd1 vssd1 vccd1 vccd1 _15368_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09354_ _15359_/Q _09354_/B _09354_/C vssd1 vssd1 vccd1 vccd1 _09362_/B sky130_fd_sc_hd__and3_1
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08305_ _08305_/A _08305_/B _08227_/B vssd1 vssd1 vccd1 vccd1 _08344_/A sky130_fd_sc_hd__or3b_2
X_09285_ _15347_/Q _09285_/B _09290_/C vssd1 vssd1 vccd1 vccd1 _09285_/Y sky130_fd_sc_hd__nand3_1
XFILLER_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08236_ _08116_/A _08236_/B vssd1 vssd1 vccd1 vccd1 _08236_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08167_ _14414_/A vssd1 vssd1 vccd1 vccd1 _14316_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_146_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08098_ _08098_/A vssd1 vssd1 vccd1 vccd1 _14782_/C sky130_fd_sc_hd__buf_2
XFILLER_109_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10060_ _10085_/C vssd1 vssd1 vccd1 vccd1 _10100_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13750_ _13750_/A vssd1 vssd1 vccd1 vccd1 _16057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10962_ _11099_/A vssd1 vssd1 vccd1 vccd1 _11085_/A sky130_fd_sc_hd__buf_2
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12701_ _12740_/A _12701_/B _12701_/C vssd1 vssd1 vccd1 vccd1 _12702_/A sky130_fd_sc_hd__and3_1
XFILLER_141_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13681_ _16048_/Q _13686_/C _13526_/X vssd1 vssd1 vccd1 vccd1 _13683_/C sky130_fd_sc_hd__a21o_1
X_10893_ _10902_/A _10893_/B _10893_/C vssd1 vssd1 vccd1 vccd1 _10894_/A sky130_fd_sc_hd__and3_1
X_15420_ _15484_/CLK _15420_/D vssd1 vssd1 vccd1 vccd1 _15420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12632_ _15871_/Q _12630_/C _12631_/X vssd1 vssd1 vccd1 vccd1 _12633_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15351_ _15351_/CLK _15351_/D vssd1 vssd1 vccd1 vccd1 _15351_/Q sky130_fd_sc_hd__dfxtp_2
X_12563_ _12559_/X _12560_/Y _12562_/Y _12557_/C vssd1 vssd1 vccd1 vccd1 _12565_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14302_ _14307_/A _14301_/Y _14295_/B _14296_/C vssd1 vssd1 vccd1 vccd1 _14304_/B
+ sky130_fd_sc_hd__o211a_1
X_11514_ _11515_/B _11515_/C _11515_/A vssd1 vssd1 vccd1 vccd1 _11516_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15282_ _15282_/CLK _15282_/D vssd1 vssd1 vccd1 vccd1 _15282_/Q sky130_fd_sc_hd__dfxtp_1
X_12494_ _12492_/X _12493_/Y _12488_/B _12489_/C vssd1 vssd1 vccd1 vccd1 _12496_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_144_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _11457_/C vssd1 vssd1 vccd1 vccd1 _11466_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14233_ _14227_/Y _14228_/X _14230_/B vssd1 vssd1 vccd1 vccd1 _14234_/B sky130_fd_sc_hd__o21a_1
XFILLER_109_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14164_ _14979_/A vssd1 vssd1 vccd1 vccd1 _14343_/A sky130_fd_sc_hd__clkbuf_2
X_11376_ _11382_/B _11376_/B vssd1 vssd1 vccd1 vccd1 _11378_/A sky130_fd_sc_hd__or2_1
XFILLER_125_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10327_ _15509_/Q _10391_/B _10331_/C vssd1 vssd1 vccd1 vccd1 _10327_/Y sky130_fd_sc_hd__nand3_1
X_13115_ _13115_/A vssd1 vssd1 vccd1 vccd1 _15948_/D sky130_fd_sc_hd__clkbuf_1
X_14095_ _16122_/Q _14095_/B _14099_/C vssd1 vssd1 vccd1 vccd1 _14095_/Y sky130_fd_sc_hd__nand3_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _15939_/Q _13051_/C _13099_/A vssd1 vssd1 vccd1 vccd1 _13048_/C sky130_fd_sc_hd__a21o_1
X_10258_ _10256_/Y _10251_/C _10253_/X _10254_/Y vssd1 vssd1 vccd1 vccd1 _10259_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_79_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _10210_/A _10189_/B _10189_/C vssd1 vssd1 vccd1 vccd1 _10190_/A sky130_fd_sc_hd__and3_1
XFILLER_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14997_ hold33/X _14997_/B vssd1 vssd1 vccd1 vccd1 _14998_/B sky130_fd_sc_hd__nor2_1
X_13948_ _13942_/B _13943_/C _13952_/A _13946_/Y vssd1 vssd1 vccd1 vccd1 _13952_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13879_ _16085_/Q _13885_/C _14587_/B vssd1 vssd1 vccd1 vccd1 _13881_/C sky130_fd_sc_hd__a21o_1
X_15618_ _15194_/Q _15618_/D vssd1 vssd1 vccd1 vccd1 _15618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15549_ _15655_/CLK _15549_/D vssd1 vssd1 vccd1 vccd1 _15549_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_148_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ _09070_/A _09070_/B vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__nor2_1
XFILLER_148_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ _08021_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08041_/A sky130_fd_sc_hd__xor2_4
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09972_ _15455_/Q _10029_/B _09979_/C vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__and3_1
XFILLER_130_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08923_ _08916_/B _08917_/C _08919_/X _08921_/Y vssd1 vssd1 vccd1 vccd1 _08924_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_97_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08854_ _15282_/Q _08859_/C _08616_/X vssd1 vssd1 vccd1 vccd1 _08856_/C sky130_fd_sc_hd__a21o_1
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07805_ _14380_/C _08027_/B vssd1 vssd1 vccd1 vccd1 _07807_/B sky130_fd_sc_hd__xnor2_1
X_08785_ _08821_/A _08785_/B _08785_/C vssd1 vssd1 vccd1 vccd1 _08786_/A sky130_fd_sc_hd__and3_1
XFILLER_85_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07736_ _07737_/A _07738_/B vssd1 vssd1 vccd1 vccd1 _07739_/A sky130_fd_sc_hd__or2_2
XFILLER_26_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07667_ _07667_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07668_/B sky130_fd_sc_hd__nor2_1
XFILLER_111_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09406_ _15365_/Q _09524_/B _09411_/C vssd1 vssd1 vccd1 vccd1 _09406_/Y sky130_fd_sc_hd__nand3_1
XFILLER_41_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07598_ _13930_/A vssd1 vssd1 vccd1 vccd1 _14459_/A sky130_fd_sc_hd__buf_2
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09337_ _09345_/A _09337_/B _09337_/C vssd1 vssd1 vccd1 vccd1 _09338_/A sky130_fd_sc_hd__and3_1
XFILLER_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09268_ _09268_/A vssd1 vssd1 vccd1 vccd1 _15344_/D sky130_fd_sc_hd__clkbuf_1
X_08219_ _08219_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08220_/B sky130_fd_sc_hd__xor2_2
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ _09236_/C vssd1 vssd1 vccd1 vccd1 _09242_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ _12377_/A vssd1 vssd1 vccd1 vccd1 _11230_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11161_ _15640_/Q _11161_/B _11169_/C vssd1 vssd1 vccd1 vccd1 _11166_/A sky130_fd_sc_hd__and3_1
XFILLER_134_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10112_ _10338_/A _10115_/C vssd1 vssd1 vccd1 vccd1 _10112_/X sky130_fd_sc_hd__or2_1
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11092_ _11090_/A _11090_/B _11091_/X vssd1 vssd1 vccd1 vccd1 _15627_/D sky130_fd_sc_hd__a21oi_1
XFILLER_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10043_ _15466_/Q _10220_/B _10043_/C vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__and3_1
X_14920_ _14920_/A _14920_/B vssd1 vssd1 vccd1 vccd1 _14921_/B sky130_fd_sc_hd__nor2_1
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14851_ _14851_/A _14851_/B vssd1 vssd1 vccd1 vccd1 _16284_/D sky130_fd_sc_hd__nor2_1
X_13802_ _13808_/A _13800_/Y _13801_/Y _13797_/C vssd1 vssd1 vccd1 vccd1 _13804_/B
+ sky130_fd_sc_hd__o211a_1
X_14782_ hold12/A _14941_/B _14782_/C vssd1 vssd1 vccd1 vccd1 _14785_/B sky130_fd_sc_hd__nand3_1
XFILLER_56_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11994_ _15769_/Q _12223_/B _12000_/C vssd1 vssd1 vccd1 vccd1 _11994_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13733_ _13734_/B _13734_/C _13734_/A vssd1 vssd1 vccd1 vccd1 _13735_/B sky130_fd_sc_hd__a21o_1
XFILLER_90_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10945_ _10945_/A vssd1 vssd1 vccd1 vccd1 _15605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13664_ _13664_/A _13664_/B _13664_/C vssd1 vssd1 vccd1 vccd1 _13665_/A sky130_fd_sc_hd__and3_1
XFILLER_32_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10876_ _15596_/Q _10876_/B _10882_/C vssd1 vssd1 vccd1 vccd1 _10879_/B sky130_fd_sc_hd__nand3_1
X_15403_ _15484_/CLK _15403_/D vssd1 vssd1 vccd1 vccd1 _15403_/Q sky130_fd_sc_hd__dfxtp_1
X_12615_ _15869_/Q _12675_/B _12623_/C vssd1 vssd1 vccd1 vccd1 _12615_/X sky130_fd_sc_hd__and3_1
X_13595_ _13595_/A _13595_/B _13595_/C vssd1 vssd1 vccd1 vccd1 _13596_/A sky130_fd_sc_hd__and3_1
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _15337_/CLK _15334_/D vssd1 vssd1 vccd1 vccd1 _15334_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12546_ _15858_/Q _12720_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12546_/X sky130_fd_sc_hd__and3_1
XFILLER_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15265_ _15274_/CLK _15265_/D vssd1 vssd1 vccd1 vccd1 _15265_/Q sky130_fd_sc_hd__dfxtp_1
X_12477_ _15845_/Q vssd1 vssd1 vccd1 vccd1 _12492_/C sky130_fd_sc_hd__inv_2
XANTENNA_4 state1[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _16149_/Q _14256_/B _14216_/C vssd1 vssd1 vccd1 vccd1 _14223_/A sky130_fd_sc_hd__and3_1
X_11428_ _11434_/A _11426_/Y _11427_/Y _11420_/C vssd1 vssd1 vccd1 vccd1 _11430_/B
+ sky130_fd_sc_hd__o211a_1
X_15196_ _15195_/Q _15196_/D vssd1 vssd1 vccd1 vccd1 _15196_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11359_ _11359_/A vssd1 vssd1 vccd1 vccd1 _15669_/D sky130_fd_sc_hd__clkbuf_1
X_14147_ _13912_/X _14145_/B _14146_/Y vssd1 vssd1 vccd1 vccd1 _16131_/D sky130_fd_sc_hd__o21a_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14078_ _14123_/A _14078_/B _14078_/C vssd1 vssd1 vccd1 vccd1 _14079_/A sky130_fd_sc_hd__and3_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _13029_/A vssd1 vssd1 vccd1 vccd1 _13283_/A sky130_fd_sc_hd__buf_2
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08570_ _08568_/Y _08564_/C _08566_/X _08567_/Y vssd1 vssd1 vccd1 vccd1 _08571_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09122_ _09120_/Y _09115_/C _09128_/A _09119_/Y vssd1 vssd1 vccd1 vccd1 _09128_/B
+ sky130_fd_sc_hd__a211oi_1
X_09053_ _15312_/Q _09061_/C _08873_/X vssd1 vssd1 vccd1 vccd1 _09053_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08004_ _13162_/C _07843_/B _07842_/A vssd1 vssd1 vccd1 vccd1 _08010_/A sky130_fd_sc_hd__o21a_1
XFILLER_129_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09955_ _09955_/A _09955_/B _09955_/C vssd1 vssd1 vccd1 vccd1 _09956_/C sky130_fd_sc_hd__nand3_1
XFILLER_106_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08906_ _08945_/C vssd1 vssd1 vccd1 vccd1 _08951_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_106_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09922_/A _09886_/B _09886_/C vssd1 vssd1 vccd1 vccd1 _09887_/A sky130_fd_sc_hd__and3_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _08835_/A _08835_/B _08836_/X vssd1 vssd1 vccd1 vccd1 _15277_/D sky130_fd_sc_hd__a21oi_1
XFILLER_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08768_ _09924_/A vssd1 vssd1 vccd1 vccd1 _09001_/B sky130_fd_sc_hd__clkbuf_2
X_07719_ _15288_/Q vssd1 vssd1 vccd1 vccd1 _08966_/A sky130_fd_sc_hd__inv_2
XFILLER_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08699_ _15258_/Q _08872_/B _08706_/C vssd1 vssd1 vccd1 vccd1 _08699_/X sky130_fd_sc_hd__and3_1
XFILLER_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10730_ _10727_/X _10728_/Y _10729_/Y _10725_/C vssd1 vssd1 vccd1 vccd1 _10732_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10661_ _11582_/A vssd1 vssd1 vccd1 vccd1 _10888_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12400_ _15834_/Q _12405_/C _12285_/X vssd1 vssd1 vccd1 vccd1 _12400_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13380_ _15995_/Q _13484_/B _13380_/C vssd1 vssd1 vccd1 vccd1 _13380_/X sky130_fd_sc_hd__and3_1
X_10592_ _10593_/B _10593_/C _10593_/A vssd1 vssd1 vccd1 vccd1 _10594_/B sky130_fd_sc_hd__a21o_1
XFILLER_127_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12331_ _15824_/Q _12391_/B _12339_/C vssd1 vssd1 vccd1 vccd1 _12331_/X sky130_fd_sc_hd__and3_1
X_12262_ _15813_/Q _12434_/B _12262_/C vssd1 vssd1 vccd1 vccd1 _12262_/X sky130_fd_sc_hd__and3_1
X_15050_ _15050_/A vssd1 vssd1 vccd1 vccd1 _15189_/B sky130_fd_sc_hd__clkbuf_2
X_11213_ _11213_/A vssd1 vssd1 vccd1 vccd1 _11228_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14001_ _13999_/A _13999_/B _13998_/Y _14000_/Y vssd1 vssd1 vccd1 vccd1 _16102_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ _12193_/A vssd1 vssd1 vccd1 vccd1 _12208_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11144_ _15637_/Q _11143_/C _10911_/X vssd1 vssd1 vccd1 vccd1 _11145_/B sky130_fd_sc_hd__a21oi_1
XFILLER_122_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11075_ _11073_/Y _11069_/C _11071_/X _11072_/Y vssd1 vssd1 vccd1 vccd1 _11076_/C
+ sky130_fd_sc_hd__a211o_1
X_15952_ _16119_/CLK _15952_/D vssd1 vssd1 vccd1 vccd1 _15952_/Q sky130_fd_sc_hd__dfxtp_1
X_10026_ _10024_/Y _10020_/C _10022_/X _10023_/Y vssd1 vssd1 vccd1 vccd1 _10027_/C
+ sky130_fd_sc_hd__a211o_1
X_14903_ _16301_/Q _14977_/B _14905_/C vssd1 vssd1 vccd1 vccd1 _14908_/A sky130_fd_sc_hd__and3_1
XFILLER_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15883_ _07603_/A _15883_/D vssd1 vssd1 vccd1 vccd1 _15883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14834_ _16285_/Q _14838_/C _14789_/X vssd1 vssd1 vccd1 vccd1 _14834_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14765_ _14765_/A _14769_/C vssd1 vssd1 vccd1 vccd1 _14768_/A sky130_fd_sc_hd__and2_1
X_11977_ _11977_/A vssd1 vssd1 vccd1 vccd1 _15766_/D sky130_fd_sc_hd__clkbuf_1
X_13716_ _14106_/A _13716_/B _13716_/C vssd1 vssd1 vccd1 vccd1 _13718_/B sky130_fd_sc_hd__or3_1
XFILLER_31_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10928_ _10963_/B vssd1 vssd1 vccd1 vccd1 _10970_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14696_ _14694_/X _14691_/A _14695_/X vssd1 vssd1 vccd1 vccd1 _14697_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13647_ _13647_/A vssd1 vssd1 vccd1 vccd1 _16039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10859_ _10859_/A _10859_/B vssd1 vssd1 vccd1 vccd1 _10863_/C sky130_fd_sc_hd__nor2_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16367_/CLK _16366_/D vssd1 vssd1 vccd1 vccd1 _16366_/Q sky130_fd_sc_hd__dfxtp_1
X_13578_ _16030_/Q _13583_/C _13526_/X vssd1 vssd1 vccd1 vccd1 _13580_/C sky130_fd_sc_hd__a21o_1
XFILLER_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15317_ _16317_/CLK _15317_/D vssd1 vssd1 vccd1 vccd1 _15317_/Q sky130_fd_sc_hd__dfxtp_1
X_12529_ _12565_/A _12529_/B _12529_/C vssd1 vssd1 vccd1 vccd1 _12530_/A sky130_fd_sc_hd__and3_1
X_16297_ _16312_/CLK _16297_/D vssd1 vssd1 vccd1 vccd1 _16297_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15248_ _15351_/CLK _15248_/D vssd1 vssd1 vccd1 vccd1 _15248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _15179_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15180_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09740_ _15419_/Q _09740_/B _09748_/C vssd1 vssd1 vccd1 vccd1 _09740_/X sky130_fd_sc_hd__and3_1
XFILLER_140_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
.ends

