VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO snn
  CLASS BLOCK ;
  FOREIGN snn ;
  ORIGIN 0.000 0.000 ;
  SIZE 419.325 BY 430.045 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.325 254.740 419.325 255.940 ;
    END
  END clk
  PIN in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 0.000 109.990 4.000 ;
    END
  END in1[0]
  PIN in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.940 4.000 351.140 ;
    END
  END in1[1]
  PIN in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.540 4.000 58.740 ;
    END
  END in1[2]
  PIN in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.610 0.000 332.170 4.000 ;
    END
  END in1[3]
  PIN in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.140 4.000 174.340 ;
    END
  END in1[4]
  PIN in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.340 4.000 116.540 ;
    END
  END in1[5]
  PIN in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.325 139.140 419.325 140.340 ;
    END
  END in1[6]
  PIN in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 426.045 142.190 430.045 ;
    END
  END in1[7]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.810 426.045 364.370 430.045 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.550 426.045 419.110 430.045 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.070 426.045 309.630 430.045 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.325 20.140 419.325 21.340 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.870 0.000 277.430 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 426.045 32.710 430.045 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.350 0.000 386.910 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.330 426.045 254.890 430.045 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 0.000 55.250 4.000 ;
    END
  END io_oeb[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.890 426.045 87.450 430.045 ;
    END
  END reset
  PIN spike_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.325 77.940 419.325 79.140 ;
    END
  END spike_out[0]
  PIN spike_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 0.000 164.730 4.000 ;
    END
  END spike_out[1]
  PIN state1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.325 312.540 419.325 313.740 ;
    END
  END state1[0]
  PIN state1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.325 370.340 419.325 371.540 ;
    END
  END state1[1]
  PIN state1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.740 4.000 289.940 ;
    END
  END state1[2]
  PIN state1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 426.045 200.150 430.045 ;
    END
  END state1[3]
  PIN state1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 0.000 219.470 4.000 ;
    END
  END state1[4]
  PIN state1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.940 4.000 232.140 ;
    END
  END state1[5]
  PIN state1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.740 4.000 408.940 ;
    END
  END state1[6]
  PIN state1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.325 196.940 419.325 198.140 ;
    END
  END state1[7]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 419.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 419.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 419.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 419.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 419.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 419.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 413.540 418.965 ;
      LAYER met1 ;
        RECT 0.070 10.640 418.990 419.120 ;
      LAYER met2 ;
        RECT 0.100 425.765 31.870 426.770 ;
        RECT 32.990 425.765 86.610 426.770 ;
        RECT 87.730 425.765 141.350 426.770 ;
        RECT 142.470 425.765 199.310 426.770 ;
        RECT 200.430 425.765 254.050 426.770 ;
        RECT 255.170 425.765 308.790 426.770 ;
        RECT 309.910 425.765 363.530 426.770 ;
        RECT 364.650 425.765 418.270 426.770 ;
        RECT 0.100 4.280 418.960 425.765 ;
        RECT 0.790 4.000 54.410 4.280 ;
        RECT 55.530 4.000 109.150 4.280 ;
        RECT 110.270 4.000 163.890 4.280 ;
        RECT 165.010 4.000 218.630 4.280 ;
        RECT 219.750 4.000 276.590 4.280 ;
        RECT 277.710 4.000 331.330 4.280 ;
        RECT 332.450 4.000 386.070 4.280 ;
        RECT 387.190 4.000 418.960 4.280 ;
      LAYER met3 ;
        RECT 4.000 409.340 415.325 419.045 ;
        RECT 4.400 407.340 415.325 409.340 ;
        RECT 4.000 371.940 415.325 407.340 ;
        RECT 4.000 369.940 414.925 371.940 ;
        RECT 4.000 351.540 415.325 369.940 ;
        RECT 4.400 349.540 415.325 351.540 ;
        RECT 4.000 314.140 415.325 349.540 ;
        RECT 4.000 312.140 414.925 314.140 ;
        RECT 4.000 290.340 415.325 312.140 ;
        RECT 4.400 288.340 415.325 290.340 ;
        RECT 4.000 256.340 415.325 288.340 ;
        RECT 4.000 254.340 414.925 256.340 ;
        RECT 4.000 232.540 415.325 254.340 ;
        RECT 4.400 230.540 415.325 232.540 ;
        RECT 4.000 198.540 415.325 230.540 ;
        RECT 4.000 196.540 414.925 198.540 ;
        RECT 4.000 174.740 415.325 196.540 ;
        RECT 4.400 172.740 415.325 174.740 ;
        RECT 4.000 140.740 415.325 172.740 ;
        RECT 4.000 138.740 414.925 140.740 ;
        RECT 4.000 116.940 415.325 138.740 ;
        RECT 4.400 114.940 415.325 116.940 ;
        RECT 4.000 79.540 415.325 114.940 ;
        RECT 4.000 77.540 414.925 79.540 ;
        RECT 4.000 59.140 415.325 77.540 ;
        RECT 4.400 57.140 415.325 59.140 ;
        RECT 4.000 21.740 415.325 57.140 ;
        RECT 4.000 19.740 414.925 21.740 ;
        RECT 4.000 10.715 415.325 19.740 ;
      LAYER met4 ;
        RECT 47.215 55.255 97.440 413.945 ;
        RECT 99.840 55.255 174.240 413.945 ;
        RECT 176.640 55.255 251.040 413.945 ;
        RECT 253.440 55.255 327.840 413.945 ;
        RECT 330.240 55.255 388.865 413.945 ;
  END
END snn
END LIBRARY

