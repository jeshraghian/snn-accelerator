magic
tech sky130A
magscale 1 2
timestamp 1654693729
<< obsli1 >>
rect 1104 2159 82708 83793
<< obsm1 >>
rect 14 2128 83798 83824
<< metal2 >>
rect 6430 85209 6542 86009
rect 17378 85209 17490 86009
rect 28326 85209 28438 86009
rect 39918 85209 40030 86009
rect 50866 85209 50978 86009
rect 61814 85209 61926 86009
rect 72762 85209 72874 86009
rect 83710 85209 83822 86009
rect -10 0 102 800
rect 10938 0 11050 800
rect 21886 0 21998 800
rect 32834 0 32946 800
rect 43782 0 43894 800
rect 55374 0 55486 800
rect 66322 0 66434 800
rect 77270 0 77382 800
<< obsm2 >>
rect 20 85153 6374 85354
rect 6598 85153 17322 85354
rect 17546 85153 28270 85354
rect 28494 85153 39862 85354
rect 40086 85153 50810 85354
rect 51034 85153 61758 85354
rect 61982 85153 72706 85354
rect 72930 85153 83654 85354
rect 20 856 83792 85153
rect 158 800 10882 856
rect 11106 800 21830 856
rect 22054 800 32778 856
rect 33002 800 43726 856
rect 43950 800 55318 856
rect 55542 800 66266 856
rect 66490 800 77214 856
rect 77438 800 83792 856
<< metal3 >>
rect 0 81548 800 81788
rect 83065 74068 83865 74308
rect 0 69988 800 70228
rect 83065 62508 83865 62748
rect 0 57748 800 57988
rect 83065 50948 83865 51188
rect 0 46188 800 46428
rect 83065 39388 83865 39628
rect 0 34628 800 34868
rect 83065 27828 83865 28068
rect 0 23068 800 23308
rect 83065 15588 83865 15828
rect 0 11508 800 11748
rect 83065 4028 83865 4268
<< obsm3 >>
rect 800 81868 83065 83809
rect 880 81468 83065 81868
rect 800 74388 83065 81468
rect 800 73988 82985 74388
rect 800 70308 83065 73988
rect 880 69908 83065 70308
rect 800 62828 83065 69908
rect 800 62428 82985 62828
rect 800 58068 83065 62428
rect 880 57668 83065 58068
rect 800 51268 83065 57668
rect 800 50868 82985 51268
rect 800 46508 83065 50868
rect 880 46108 83065 46508
rect 800 39708 83065 46108
rect 800 39308 82985 39708
rect 800 34948 83065 39308
rect 880 34548 83065 34948
rect 800 28148 83065 34548
rect 800 27748 82985 28148
rect 800 23388 83065 27748
rect 880 22988 83065 23388
rect 800 15908 83065 22988
rect 800 15508 82985 15908
rect 800 11828 83065 15508
rect 880 11428 83065 11828
rect 800 4348 83065 11428
rect 800 3948 82985 4348
rect 800 2143 83065 3948
<< metal4 >>
rect 4208 2128 4528 83824
rect 19568 2128 19888 83824
rect 34928 2128 35248 83824
rect 50288 2128 50608 83824
rect 65648 2128 65968 83824
rect 81008 2128 81328 83824
<< obsm4 >>
rect 9443 11051 19488 82789
rect 19968 11051 34848 82789
rect 35328 11051 50208 82789
rect 50688 11051 65568 82789
rect 66048 11051 77773 82789
<< labels >>
rlabel metal3 s 83065 50948 83865 51188 6 clk
port 1 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 in1[0]
port 2 nsew signal input
rlabel metal3 s 0 69988 800 70228 6 in1[1]
port 3 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 in1[2]
port 4 nsew signal input
rlabel metal2 s 66322 0 66434 800 6 in1[3]
port 5 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 in1[4]
port 6 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 in1[5]
port 7 nsew signal input
rlabel metal3 s 83065 27828 83865 28068 6 in1[6]
port 8 nsew signal input
rlabel metal2 s 28326 85209 28438 86009 6 in1[7]
port 9 nsew signal input
rlabel metal2 s -10 0 102 800 6 io_oeb[0]
port 10 nsew signal output
rlabel metal2 s 72762 85209 72874 86009 6 io_oeb[1]
port 11 nsew signal output
rlabel metal2 s 83710 85209 83822 86009 6 io_oeb[2]
port 12 nsew signal output
rlabel metal2 s 61814 85209 61926 86009 6 io_oeb[3]
port 13 nsew signal output
rlabel metal3 s 83065 4028 83865 4268 6 io_oeb[4]
port 14 nsew signal output
rlabel metal2 s 55374 0 55486 800 6 io_oeb[5]
port 15 nsew signal output
rlabel metal2 s 6430 85209 6542 86009 6 io_oeb[6]
port 16 nsew signal output
rlabel metal2 s 77270 0 77382 800 6 io_oeb[7]
port 17 nsew signal output
rlabel metal2 s 50866 85209 50978 86009 6 io_oeb[8]
port 18 nsew signal output
rlabel metal2 s 10938 0 11050 800 6 io_oeb[9]
port 19 nsew signal output
rlabel metal2 s 17378 85209 17490 86009 6 reset
port 20 nsew signal input
rlabel metal3 s 83065 15588 83865 15828 6 spike_out[0]
port 21 nsew signal output
rlabel metal2 s 32834 0 32946 800 6 spike_out[1]
port 22 nsew signal output
rlabel metal3 s 83065 62508 83865 62748 6 state1[0]
port 23 nsew signal output
rlabel metal3 s 83065 74068 83865 74308 6 state1[1]
port 24 nsew signal output
rlabel metal3 s 0 57748 800 57988 6 state1[2]
port 25 nsew signal output
rlabel metal2 s 39918 85209 40030 86009 6 state1[3]
port 26 nsew signal output
rlabel metal2 s 43782 0 43894 800 6 state1[4]
port 27 nsew signal output
rlabel metal3 s 0 46188 800 46428 6 state1[5]
port 28 nsew signal output
rlabel metal3 s 0 81548 800 81788 6 state1[6]
port 29 nsew signal output
rlabel metal3 s 83065 39388 83865 39628 6 state1[7]
port 30 nsew signal output
rlabel metal4 s 4208 2128 4528 83824 6 vccd1
port 31 nsew power input
rlabel metal4 s 34928 2128 35248 83824 6 vccd1
port 31 nsew power input
rlabel metal4 s 65648 2128 65968 83824 6 vccd1
port 31 nsew power input
rlabel metal4 s 19568 2128 19888 83824 6 vssd1
port 32 nsew ground input
rlabel metal4 s 50288 2128 50608 83824 6 vssd1
port 32 nsew ground input
rlabel metal4 s 81008 2128 81328 83824 6 vssd1
port 32 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 83865 86009
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 22963898
string GDS_FILE /openlane/designs/snn/runs/RUN_2022.06.08_12.57.24/results/finishing/snn.magic.gds
string GDS_START 563548
<< end >>

