VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_snn
  CLASS BLOCK ;
  FOREIGN wrapped_snn ;
  ORIGIN 0.000 0.000 ;
  SIZE 422.705 BY 433.425 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 417.940 422.705 419.140 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 98.340 422.705 99.540 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 429.425 48.810 433.425 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.140 4.000 242.340 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.910 429.425 380.470 433.425 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.070 429.425 309.630 433.425 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.740 4.000 272.940 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.540 4.000 75.740 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 429.425 148.630 433.425 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 0.000 113.210 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.540 4.000 58.740 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 387.340 422.705 388.540 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 6.540 422.705 7.740 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.030 429.425 367.590 433.425 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.340 4.000 303.540 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.140 4.000 395.340 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 190.140 422.705 191.340 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.940 4.000 45.140 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.140 4.000 412.340 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 429.425 206.590 433.425 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 404.340 422.705 405.540 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.450 0.000 403.010 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 128.940 422.705 130.140 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 429.425 193.710 433.425 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.550 0.000 258.110 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 220.740 422.705 221.940 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.140 4.000 259.340 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.770 0.000 100.330 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.730 0.000 158.290 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 37.140 422.705 38.340 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.940 4.000 334.140 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 429.425 135.750 433.425 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 142.540 422.705 143.740 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 234.340 422.705 235.540 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.010 429.425 235.570 433.425 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 173.140 422.705 174.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.110 429.425 251.670 433.425 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 429.425 280.650 433.425 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.050 429.425 338.610 433.425 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.770 429.425 422.330 433.425 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 356.740 422.705 357.940 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 0.000 55.250 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 429.425 77.790 433.425 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 0.000 187.270 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 0.000 245.230 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 373.740 422.705 374.940 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.470 0.000 374.030 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 281.940 422.705 283.140 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.050 429.425 177.610 433.425 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.540 4.000 211.740 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 429.425 106.770 433.425 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.130 429.425 222.690 433.425 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.610 0.000 332.170 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 0.000 129.310 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 111.940 422.705 113.140 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 429.425 119.650 433.425 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 295.540 422.705 296.740 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 0.000 26.270 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.570 0.000 390.130 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 81.340 422.705 82.540 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.890 429.425 409.450 433.425 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.540 4.000 364.740 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.490 0.000 345.050 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 0.000 171.170 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.940 4.000 351.140 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 326.140 422.705 327.340 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.940 4.000 198.140 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 20.140 422.705 21.340 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 429.425 6.950 433.425 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 429.425 61.690 433.425 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.740 4.000 289.940 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.630 0.000 303.190 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 0.000 42.370 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.940 4.000 181.140 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.550 0.000 419.110 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 251.340 422.705 252.540 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 159.540 422.705 160.740 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.510 0.000 316.070 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.340 4.000 320.540 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 67.740 422.705 68.940 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.540 4.000 228.740 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 312.540 422.705 313.740 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.590 0.000 361.150 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 343.140 422.705 344.340 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.690 0.000 216.250 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.140 4.000 89.340 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.340 4.000 167.540 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.650 0.000 274.210 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 429.425 32.710 433.425 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 429.425 164.730 433.425 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.970 429.425 293.530 433.425 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.940 4.000 28.140 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 0.000 71.350 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 0.000 13.390 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.930 429.425 351.490 433.425 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 429.425 264.550 433.425 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 0.000 200.150 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.010 429.425 396.570 433.425 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 50.740 422.705 51.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.740 4.000 425.940 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.340 4.000 150.540 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 0.000 84.230 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 0.000 142.190 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.740 4.000 136.940 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 264.940 422.705 266.140 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 0.000 229.130 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.140 4.000 106.340 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.950 429.425 322.510 433.425 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 429.425 19.830 433.425 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 429.425 90.670 433.425 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.530 0.000 287.090 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.740 4.000 119.940 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.540 4.000 381.740 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 421.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 421.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 421.840 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 421.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 421.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 421.840 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 418.705 203.740 422.705 204.940 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 416.760 421.685 ;
      LAYER met1 ;
        RECT 0.070 9.560 422.210 421.840 ;
      LAYER met2 ;
        RECT 0.100 429.145 6.110 430.170 ;
        RECT 7.230 429.145 18.990 430.170 ;
        RECT 20.110 429.145 31.870 430.170 ;
        RECT 32.990 429.145 47.970 430.170 ;
        RECT 49.090 429.145 60.850 430.170 ;
        RECT 61.970 429.145 76.950 430.170 ;
        RECT 78.070 429.145 89.830 430.170 ;
        RECT 90.950 429.145 105.930 430.170 ;
        RECT 107.050 429.145 118.810 430.170 ;
        RECT 119.930 429.145 134.910 430.170 ;
        RECT 136.030 429.145 147.790 430.170 ;
        RECT 148.910 429.145 163.890 430.170 ;
        RECT 165.010 429.145 176.770 430.170 ;
        RECT 177.890 429.145 192.870 430.170 ;
        RECT 193.990 429.145 205.750 430.170 ;
        RECT 206.870 429.145 221.850 430.170 ;
        RECT 222.970 429.145 234.730 430.170 ;
        RECT 235.850 429.145 250.830 430.170 ;
        RECT 251.950 429.145 263.710 430.170 ;
        RECT 264.830 429.145 279.810 430.170 ;
        RECT 280.930 429.145 292.690 430.170 ;
        RECT 293.810 429.145 308.790 430.170 ;
        RECT 309.910 429.145 321.670 430.170 ;
        RECT 322.790 429.145 337.770 430.170 ;
        RECT 338.890 429.145 350.650 430.170 ;
        RECT 351.770 429.145 366.750 430.170 ;
        RECT 367.870 429.145 379.630 430.170 ;
        RECT 380.750 429.145 395.730 430.170 ;
        RECT 396.850 429.145 408.610 430.170 ;
        RECT 409.730 429.145 421.490 430.170 ;
        RECT 0.100 4.280 422.180 429.145 ;
        RECT 0.790 4.000 12.550 4.280 ;
        RECT 13.670 4.000 25.430 4.280 ;
        RECT 26.550 4.000 41.530 4.280 ;
        RECT 42.650 4.000 54.410 4.280 ;
        RECT 55.530 4.000 70.510 4.280 ;
        RECT 71.630 4.000 83.390 4.280 ;
        RECT 84.510 4.000 99.490 4.280 ;
        RECT 100.610 4.000 112.370 4.280 ;
        RECT 113.490 4.000 128.470 4.280 ;
        RECT 129.590 4.000 141.350 4.280 ;
        RECT 142.470 4.000 157.450 4.280 ;
        RECT 158.570 4.000 170.330 4.280 ;
        RECT 171.450 4.000 186.430 4.280 ;
        RECT 187.550 4.000 199.310 4.280 ;
        RECT 200.430 4.000 215.410 4.280 ;
        RECT 216.530 4.000 228.290 4.280 ;
        RECT 229.410 4.000 244.390 4.280 ;
        RECT 245.510 4.000 257.270 4.280 ;
        RECT 258.390 4.000 273.370 4.280 ;
        RECT 274.490 4.000 286.250 4.280 ;
        RECT 287.370 4.000 302.350 4.280 ;
        RECT 303.470 4.000 315.230 4.280 ;
        RECT 316.350 4.000 331.330 4.280 ;
        RECT 332.450 4.000 344.210 4.280 ;
        RECT 345.330 4.000 360.310 4.280 ;
        RECT 361.430 4.000 373.190 4.280 ;
        RECT 374.310 4.000 389.290 4.280 ;
        RECT 390.410 4.000 402.170 4.280 ;
        RECT 403.290 4.000 418.270 4.280 ;
        RECT 419.390 4.000 422.180 4.280 ;
      LAYER met3 ;
        RECT 4.400 424.340 418.705 425.505 ;
        RECT 4.000 419.540 418.705 424.340 ;
        RECT 4.000 417.540 418.305 419.540 ;
        RECT 4.000 412.740 418.705 417.540 ;
        RECT 4.400 410.740 418.705 412.740 ;
        RECT 4.000 405.940 418.705 410.740 ;
        RECT 4.000 403.940 418.305 405.940 ;
        RECT 4.000 395.740 418.705 403.940 ;
        RECT 4.400 393.740 418.705 395.740 ;
        RECT 4.000 388.940 418.705 393.740 ;
        RECT 4.000 386.940 418.305 388.940 ;
        RECT 4.000 382.140 418.705 386.940 ;
        RECT 4.400 380.140 418.705 382.140 ;
        RECT 4.000 375.340 418.705 380.140 ;
        RECT 4.000 373.340 418.305 375.340 ;
        RECT 4.000 365.140 418.705 373.340 ;
        RECT 4.400 363.140 418.705 365.140 ;
        RECT 4.000 358.340 418.705 363.140 ;
        RECT 4.000 356.340 418.305 358.340 ;
        RECT 4.000 351.540 418.705 356.340 ;
        RECT 4.400 349.540 418.705 351.540 ;
        RECT 4.000 344.740 418.705 349.540 ;
        RECT 4.000 342.740 418.305 344.740 ;
        RECT 4.000 334.540 418.705 342.740 ;
        RECT 4.400 332.540 418.705 334.540 ;
        RECT 4.000 327.740 418.705 332.540 ;
        RECT 4.000 325.740 418.305 327.740 ;
        RECT 4.000 320.940 418.705 325.740 ;
        RECT 4.400 318.940 418.705 320.940 ;
        RECT 4.000 314.140 418.705 318.940 ;
        RECT 4.000 312.140 418.305 314.140 ;
        RECT 4.000 303.940 418.705 312.140 ;
        RECT 4.400 301.940 418.705 303.940 ;
        RECT 4.000 297.140 418.705 301.940 ;
        RECT 4.000 295.140 418.305 297.140 ;
        RECT 4.000 290.340 418.705 295.140 ;
        RECT 4.400 288.340 418.705 290.340 ;
        RECT 4.000 283.540 418.705 288.340 ;
        RECT 4.000 281.540 418.305 283.540 ;
        RECT 4.000 273.340 418.705 281.540 ;
        RECT 4.400 271.340 418.705 273.340 ;
        RECT 4.000 266.540 418.705 271.340 ;
        RECT 4.000 264.540 418.305 266.540 ;
        RECT 4.000 259.740 418.705 264.540 ;
        RECT 4.400 257.740 418.705 259.740 ;
        RECT 4.000 252.940 418.705 257.740 ;
        RECT 4.000 250.940 418.305 252.940 ;
        RECT 4.000 242.740 418.705 250.940 ;
        RECT 4.400 240.740 418.705 242.740 ;
        RECT 4.000 235.940 418.705 240.740 ;
        RECT 4.000 233.940 418.305 235.940 ;
        RECT 4.000 229.140 418.705 233.940 ;
        RECT 4.400 227.140 418.705 229.140 ;
        RECT 4.000 222.340 418.705 227.140 ;
        RECT 4.000 220.340 418.305 222.340 ;
        RECT 4.000 212.140 418.705 220.340 ;
        RECT 4.400 210.140 418.705 212.140 ;
        RECT 4.000 205.340 418.705 210.140 ;
        RECT 4.000 203.340 418.305 205.340 ;
        RECT 4.000 198.540 418.705 203.340 ;
        RECT 4.400 196.540 418.705 198.540 ;
        RECT 4.000 191.740 418.705 196.540 ;
        RECT 4.000 189.740 418.305 191.740 ;
        RECT 4.000 181.540 418.705 189.740 ;
        RECT 4.400 179.540 418.705 181.540 ;
        RECT 4.000 174.740 418.705 179.540 ;
        RECT 4.000 172.740 418.305 174.740 ;
        RECT 4.000 167.940 418.705 172.740 ;
        RECT 4.400 165.940 418.705 167.940 ;
        RECT 4.000 161.140 418.705 165.940 ;
        RECT 4.000 159.140 418.305 161.140 ;
        RECT 4.000 150.940 418.705 159.140 ;
        RECT 4.400 148.940 418.705 150.940 ;
        RECT 4.000 144.140 418.705 148.940 ;
        RECT 4.000 142.140 418.305 144.140 ;
        RECT 4.000 137.340 418.705 142.140 ;
        RECT 4.400 135.340 418.705 137.340 ;
        RECT 4.000 130.540 418.705 135.340 ;
        RECT 4.000 128.540 418.305 130.540 ;
        RECT 4.000 120.340 418.705 128.540 ;
        RECT 4.400 118.340 418.705 120.340 ;
        RECT 4.000 113.540 418.705 118.340 ;
        RECT 4.000 111.540 418.305 113.540 ;
        RECT 4.000 106.740 418.705 111.540 ;
        RECT 4.400 104.740 418.705 106.740 ;
        RECT 4.000 99.940 418.705 104.740 ;
        RECT 4.000 97.940 418.305 99.940 ;
        RECT 4.000 89.740 418.705 97.940 ;
        RECT 4.400 87.740 418.705 89.740 ;
        RECT 4.000 82.940 418.705 87.740 ;
        RECT 4.000 80.940 418.305 82.940 ;
        RECT 4.000 76.140 418.705 80.940 ;
        RECT 4.400 74.140 418.705 76.140 ;
        RECT 4.000 69.340 418.705 74.140 ;
        RECT 4.000 67.340 418.305 69.340 ;
        RECT 4.000 59.140 418.705 67.340 ;
        RECT 4.400 57.140 418.705 59.140 ;
        RECT 4.000 52.340 418.705 57.140 ;
        RECT 4.000 50.340 418.305 52.340 ;
        RECT 4.000 45.540 418.705 50.340 ;
        RECT 4.400 43.540 418.705 45.540 ;
        RECT 4.000 38.740 418.705 43.540 ;
        RECT 4.000 36.740 418.305 38.740 ;
        RECT 4.000 28.540 418.705 36.740 ;
        RECT 4.400 26.540 418.705 28.540 ;
        RECT 4.000 21.740 418.705 26.540 ;
        RECT 4.000 19.740 418.305 21.740 ;
        RECT 4.000 14.940 418.705 19.740 ;
        RECT 4.400 12.940 418.705 14.940 ;
        RECT 4.000 10.715 418.705 12.940 ;
      LAYER met4 ;
        RECT 26.975 17.175 97.440 407.825 ;
        RECT 99.840 17.175 174.240 407.825 ;
        RECT 176.640 17.175 251.040 407.825 ;
        RECT 253.440 17.175 327.840 407.825 ;
        RECT 330.240 17.175 401.745 407.825 ;
  END
END wrapped_snn
END LIBRARY

